magic
tech sky130A
magscale 1 2
timestamp 1711995521
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
use trans_gate  x1
timestamp 1711994542
transform 1 0 -3618 0 1 2292
box 0 -2380 2272 590
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[0]
timestamp 1711994542
transform 1 0 8716 0 1 -6762
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[1]
timestamp 1711994542
transform 1 0 8656 0 1 -5782
box -1028 -388 1028 388
use sky130_fd_pr__nfet_01v8_BW73UN  XM2[0]
timestamp 1711994542
transform 1 0 11246 0 1 -6692
box -996 -340 996 340
use sky130_fd_pr__nfet_01v8_BW73UN  XM2[1]
timestamp 1711994542
transform 1 0 11374 0 1 -5760
box -996 -340 996 340
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[0]
timestamp 1711994542
transform -1 0 10856 0 -1 -933
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[1]
timestamp 1711994542
transform 1 0 12742 0 1 -401
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[0]
timestamp 1711994542
transform 1 0 18126 0 1 -1065
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1711994542
transform 1 0 17026 0 1 77
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[0]
timestamp 1711994542
transform 1 0 12742 0 1 -933
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[1]
timestamp 1711994542
transform 1 0 10856 0 1 -401
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[0]
timestamp 1711994542
transform 1 0 11686 0 1 4149
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1711994542
transform 1 0 11728 0 1 5149
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[2]
timestamp 1711994542
transform 1 0 11624 0 1 3089
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1711994542
transform 1 0 11842 0 1 2099
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1711994542
transform 1 0 3316 0 1 -419
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_697RXD  XM8
timestamp 1711994542
transform 1 0 1076 0 1 -5334
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1711994542
transform 1 0 6950 0 1 -1089
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1711994542
transform 1 0 4524 0 1 -5320
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1711994542
transform 1 0 10488 0 1 -4530
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1711994542
transform 1 0 5816 0 1 -4514
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1711994542
transform 1 0 970 0 1 -4440
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1711994542
transform 1 0 2824 0 1 -5366
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1711994542
transform 1 0 4250 0 1 -1353
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1711994542
transform 1 0 2840 0 1 -1417
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1711994542
transform 1 0 5716 0 1 -5382
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1711994542
transform 1 0 5426 0 1 -305
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1711994542
transform 1 0 2826 0 1 -4562
box -496 -310 496 310
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 dvdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vref
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vin
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 ibias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 vss
port 6 nsew
<< end >>

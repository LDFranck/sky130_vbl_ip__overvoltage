magic
tech sky130A
timestamp 1711651911
<< pwell >>
rect -364 -179 364 179
<< mvnmos >>
rect -250 -50 250 50
<< mvndiff >>
rect -279 44 -250 50
rect -279 -44 -273 44
rect -256 -44 -250 44
rect -279 -50 -250 -44
rect 250 44 279 50
rect 250 -44 256 44
rect 273 -44 279 44
rect 250 -50 279 -44
<< mvndiffc >>
rect -273 -44 -256 44
rect 256 -44 273 44
<< mvpsubdiff >>
rect -346 155 346 161
rect -346 138 -292 155
rect 292 138 346 155
rect -346 132 346 138
rect -346 107 -317 132
rect -346 -107 -340 107
rect -323 -107 -317 107
rect 317 107 346 132
rect -346 -132 -317 -107
rect 317 -107 323 107
rect 340 -107 346 107
rect 317 -132 346 -107
rect -346 -138 346 -132
rect -346 -155 -292 -138
rect 292 -155 346 -138
rect -346 -161 346 -155
<< mvpsubdiffcont >>
rect -292 138 292 155
rect -340 -107 -323 107
rect 323 -107 340 107
rect -292 -155 292 -138
<< poly >>
rect -250 86 250 94
rect -250 69 -242 86
rect 242 69 250 86
rect -250 50 250 69
rect -250 -69 250 -50
rect -250 -86 -242 -69
rect 242 -86 250 -69
rect -250 -94 250 -86
<< polycont >>
rect -242 69 242 86
rect -242 -86 242 -69
<< locali >>
rect -340 138 -292 155
rect 292 138 340 155
rect -340 107 -323 138
rect 323 107 340 138
rect -250 69 -242 86
rect 242 69 250 86
rect -273 44 -256 52
rect -273 -52 -256 -44
rect 256 44 273 52
rect 256 -52 273 -44
rect -250 -86 -242 -69
rect 242 -86 250 -69
rect -340 -138 -323 -107
rect 323 -138 340 -107
rect -340 -155 -292 -138
rect 292 -155 340 -138
<< viali >>
rect -242 69 242 86
rect -273 -44 -256 44
rect 256 -44 273 44
rect -242 -86 242 -69
<< metal1 >>
rect -248 86 248 89
rect -248 69 -242 86
rect 242 69 248 86
rect -248 66 248 69
rect -276 44 -253 50
rect -276 -44 -273 44
rect -256 -44 -253 44
rect -276 -50 -253 -44
rect 253 44 276 50
rect 253 -44 256 44
rect 273 -44 276 44
rect 253 -50 276 -44
rect -248 -69 248 -66
rect -248 -86 -242 -69
rect 242 -86 248 -69
rect -248 -89 248 -86
<< properties >>
string FIXED_BBOX -331 -146 331 146
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

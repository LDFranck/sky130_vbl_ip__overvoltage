magic
tech sky130A
magscale 1 2
timestamp 1712240559
<< pwell >>
rect -2008 -1992 2008 1992
<< psubdiff >>
rect -1972 1922 -1876 1956
rect 1876 1922 1972 1956
rect -1972 1860 -1938 1922
rect 1938 1860 1972 1922
rect -1972 -1922 -1938 -1860
rect 1938 -1922 1972 -1860
rect -1972 -1956 -1876 -1922
rect 1876 -1956 1972 -1922
<< psubdiffcont >>
rect -1876 1922 1876 1956
rect -1972 -1860 -1938 1860
rect 1938 -1860 1972 1860
rect -1876 -1956 1876 -1922
<< xpolycontact >>
rect -1842 1394 -1560 1826
rect -1842 -1826 -1560 -1394
rect -1464 1394 -1182 1826
rect -1464 -1826 -1182 -1394
rect -1086 1394 -804 1826
rect -1086 -1826 -804 -1394
rect -708 1394 -426 1826
rect -708 -1826 -426 -1394
rect -330 1394 -48 1826
rect -330 -1826 -48 -1394
rect 48 1394 330 1826
rect 48 -1826 330 -1394
rect 426 1394 708 1826
rect 426 -1826 708 -1394
rect 804 1394 1086 1826
rect 804 -1826 1086 -1394
rect 1182 1394 1464 1826
rect 1182 -1826 1464 -1394
rect 1560 1394 1842 1826
rect 1560 -1826 1842 -1394
<< xpolyres >>
rect -1842 -1394 -1560 1394
rect -1464 -1394 -1182 1394
rect -1086 -1394 -804 1394
rect -708 -1394 -426 1394
rect -330 -1394 -48 1394
rect 48 -1394 330 1394
rect 426 -1394 708 1394
rect 804 -1394 1086 1394
rect 1182 -1394 1464 1394
rect 1560 -1394 1842 1394
<< locali >>
rect -1972 1922 -1876 1956
rect 1876 1922 1972 1956
rect -1972 1860 -1938 1922
rect 1938 1860 1972 1922
rect -1972 -1922 -1938 -1860
rect 1938 -1922 1972 -1860
rect -1972 -1956 -1876 -1922
rect 1876 -1956 1972 -1922
<< viali >>
rect -1826 1411 -1576 1808
rect -1448 1411 -1198 1808
rect -1070 1411 -820 1808
rect -692 1411 -442 1808
rect -314 1411 -64 1808
rect 64 1411 314 1808
rect 442 1411 692 1808
rect 820 1411 1070 1808
rect 1198 1411 1448 1808
rect 1576 1411 1826 1808
rect -1826 -1808 -1576 -1411
rect -1448 -1808 -1198 -1411
rect -1070 -1808 -820 -1411
rect -692 -1808 -442 -1411
rect -314 -1808 -64 -1411
rect 64 -1808 314 -1411
rect 442 -1808 692 -1411
rect 820 -1808 1070 -1411
rect 1198 -1808 1448 -1411
rect 1576 -1808 1826 -1411
<< metal1 >>
rect -1832 1808 -1570 1820
rect -1832 1411 -1826 1808
rect -1576 1411 -1570 1808
rect -1832 1399 -1570 1411
rect -1454 1808 -1192 1820
rect -1454 1411 -1448 1808
rect -1198 1411 -1192 1808
rect -1454 1399 -1192 1411
rect -1076 1808 -814 1820
rect -1076 1411 -1070 1808
rect -820 1411 -814 1808
rect -1076 1399 -814 1411
rect -698 1808 -436 1820
rect -698 1411 -692 1808
rect -442 1411 -436 1808
rect -698 1399 -436 1411
rect -320 1808 -58 1820
rect -320 1411 -314 1808
rect -64 1411 -58 1808
rect -320 1399 -58 1411
rect 58 1808 320 1820
rect 58 1411 64 1808
rect 314 1411 320 1808
rect 58 1399 320 1411
rect 436 1808 698 1820
rect 436 1411 442 1808
rect 692 1411 698 1808
rect 436 1399 698 1411
rect 814 1808 1076 1820
rect 814 1411 820 1808
rect 1070 1411 1076 1808
rect 814 1399 1076 1411
rect 1192 1808 1454 1820
rect 1192 1411 1198 1808
rect 1448 1411 1454 1808
rect 1192 1399 1454 1411
rect 1570 1808 1832 1820
rect 1570 1411 1576 1808
rect 1826 1411 1832 1808
rect 1570 1399 1832 1411
rect -1832 -1411 -1570 -1399
rect -1832 -1808 -1826 -1411
rect -1576 -1808 -1570 -1411
rect -1832 -1820 -1570 -1808
rect -1454 -1411 -1192 -1399
rect -1454 -1808 -1448 -1411
rect -1198 -1808 -1192 -1411
rect -1454 -1820 -1192 -1808
rect -1076 -1411 -814 -1399
rect -1076 -1808 -1070 -1411
rect -820 -1808 -814 -1411
rect -1076 -1820 -814 -1808
rect -698 -1411 -436 -1399
rect -698 -1808 -692 -1411
rect -442 -1808 -436 -1411
rect -698 -1820 -436 -1808
rect -320 -1411 -58 -1399
rect -320 -1808 -314 -1411
rect -64 -1808 -58 -1411
rect -320 -1820 -58 -1808
rect 58 -1411 320 -1399
rect 58 -1808 64 -1411
rect 314 -1808 320 -1411
rect 58 -1820 320 -1808
rect 436 -1411 698 -1399
rect 436 -1808 442 -1411
rect 692 -1808 698 -1411
rect 436 -1820 698 -1808
rect 814 -1411 1076 -1399
rect 814 -1808 820 -1411
rect 1070 -1808 1076 -1411
rect 814 -1820 1076 -1808
rect 1192 -1411 1454 -1399
rect 1192 -1808 1198 -1411
rect 1448 -1808 1454 -1411
rect 1192 -1820 1454 -1808
rect 1570 -1411 1832 -1399
rect 1570 -1808 1576 -1411
rect 1826 -1808 1832 -1411
rect 1570 -1820 1832 -1808
<< properties >>
string FIXED_BBOX -1955 -1939 1955 1939
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 14.1 m 1 nx 10 wmin 1.410 lmin 0.50 rho 2000 val 20.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713017665
<< nwell >>
rect -758 -897 758 897
<< mvpmos >>
rect -500 -600 500 600
<< mvpdiff >>
rect -558 588 -500 600
rect -558 -588 -546 588
rect -512 -588 -500 588
rect -558 -600 -500 -588
rect 500 588 558 600
rect 500 -588 512 588
rect 546 -588 558 588
rect 500 -600 558 -588
<< mvpdiffc >>
rect -546 -588 -512 588
rect 512 -588 546 588
<< mvnsubdiff >>
rect -692 819 692 831
rect -692 785 -584 819
rect 584 785 692 819
rect -692 773 692 785
rect -692 723 -634 773
rect -692 -723 -680 723
rect -646 -723 -634 723
rect 634 723 692 773
rect -692 -773 -634 -723
rect 634 -723 646 723
rect 680 -723 692 723
rect 634 -773 692 -723
rect -692 -785 692 -773
rect -692 -819 -584 -785
rect 584 -819 692 -785
rect -692 -831 692 -819
<< mvnsubdiffcont >>
rect -584 785 584 819
rect -680 -723 -646 723
rect 646 -723 680 723
rect -584 -819 584 -785
<< poly >>
rect -500 681 500 697
rect -500 647 -484 681
rect 484 647 500 681
rect -500 600 500 647
rect -500 -647 500 -600
rect -500 -681 -484 -647
rect 484 -681 500 -647
rect -500 -697 500 -681
<< polycont >>
rect -484 647 484 681
rect -484 -681 484 -647
<< locali >>
rect -680 785 -584 819
rect 584 785 680 819
rect -680 723 -646 785
rect 646 723 680 785
rect -500 647 -484 681
rect 484 647 500 681
rect -546 588 -512 604
rect -546 -604 -512 -588
rect 512 588 546 604
rect 512 -604 546 -588
rect -500 -681 -484 -647
rect 484 -681 500 -647
rect -680 -785 -646 -723
rect 646 -785 680 -723
rect -680 -819 -584 -785
rect 584 -819 680 -785
<< viali >>
rect -484 647 484 681
rect -546 -588 -512 588
rect 512 -588 546 588
rect -484 -681 484 -647
<< metal1 >>
rect -496 681 496 687
rect -496 647 -484 681
rect 484 647 496 681
rect -496 641 496 647
rect -552 588 -506 600
rect -552 -588 -546 588
rect -512 -588 -506 588
rect -552 -600 -506 -588
rect 506 588 552 600
rect 506 -588 512 588
rect 546 -588 552 588
rect 506 -600 552 -588
rect -496 -647 496 -641
rect -496 -681 -484 -647
rect 484 -681 496 -647
rect -496 -687 496 -681
<< properties >>
string FIXED_BBOX -663 -802 663 802
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 6.0 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713117387
<< locali >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 2319 -509 3279 -340
rect 7041 -369 8144 -340
rect 7041 -492 7262 -369
rect 8107 -492 8144 -369
rect 7041 -538 8144 -492
rect 7041 -1104 7224 -538
rect 7040 -1740 7224 -1226
rect 1183 -2314 2143 -1781
rect 7357 -2034 8144 -1774
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 7040 -2121 8144 -2034
rect 7040 -2244 7082 -2121
rect 8082 -2244 8144 -2121
rect 7040 -2314 8144 -2244
<< viali >>
rect 1223 -493 2106 -370
rect 7262 -492 8107 -369
rect 2357 -2286 3240 -2163
rect 7082 -2244 8082 -2121
<< metal1 >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 7224 -369 8144 -340
rect 7224 -492 7262 -369
rect 8107 -492 8144 -369
rect 7224 -538 8144 -492
rect 1183 -758 1325 -539
rect 1353 -710 1363 -658
rect 1963 -710 1973 -658
rect 2489 -670 2499 -618
rect 3099 -670 3109 -618
rect 1183 -959 1357 -758
rect 1969 -830 2494 -746
rect 1969 -887 2205 -830
rect 2345 -887 2494 -830
rect 1969 -958 2494 -887
rect 1183 -1362 1325 -959
rect 1353 -1058 1363 -1006
rect 1963 -1058 1973 -1006
rect 2489 -1167 2505 -1151
rect 3095 -1167 3105 -1151
rect 2489 -1219 2499 -1167
rect 3099 -1219 3105 -1167
rect 1353 -1314 1363 -1262
rect 1963 -1314 1973 -1262
rect 1183 -1562 1357 -1362
rect 1969 -1427 2461 -1362
rect 1969 -1484 1985 -1427
rect 2125 -1484 2461 -1427
rect 2489 -1457 2499 -1405
rect 3099 -1457 3105 -1405
rect 2489 -1473 2504 -1457
rect 3095 -1473 3105 -1457
rect 1969 -1562 2461 -1484
rect 2462 -1562 2493 -1505
rect 1353 -1662 1363 -1610
rect 1963 -1662 1973 -1610
rect 2271 -1905 2493 -1562
rect 2489 -1953 3109 -1937
rect 2489 -2005 2499 -1953
rect 3099 -2005 3109 -1953
rect 3137 -2115 3279 -718
rect 7224 -721 7346 -538
rect 7374 -673 7384 -621
rect 7984 -673 7994 -621
rect 7224 -921 7378 -721
rect 7990 -921 8144 -721
rect 7374 -1021 7384 -969
rect 7984 -1021 7991 -969
rect 8019 -1104 8144 -921
rect 7258 -1225 8144 -1104
rect 7258 -1226 8110 -1225
rect 7258 -1400 7349 -1226
rect 7377 -1352 7383 -1300
rect 7984 -1352 7994 -1300
rect 7377 -1368 7994 -1352
rect 7258 -1599 7326 -1400
rect 7378 -1599 7388 -1400
rect 7258 -1600 7377 -1599
rect 7990 -1600 8144 -1400
rect 7374 -1700 7384 -1648
rect 7985 -1700 7995 -1648
rect 7132 -1926 7142 -1848
rect 7282 -1926 7292 -1848
rect 8023 -2034 8144 -1600
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 7040 -2121 8144 -2034
rect 7040 -2244 7082 -2121
rect 8082 -2244 8144 -2121
rect 7040 -2313 8144 -2244
rect 7040 -2314 7357 -2313
<< via1 >>
rect 1363 -710 1963 -658
rect 2499 -670 3099 -618
rect 2205 -887 2345 -830
rect 1363 -1058 1963 -1006
rect 2499 -1219 3099 -1167
rect 1363 -1314 1963 -1262
rect 1985 -1484 2125 -1427
rect 2499 -1457 3099 -1405
rect 1363 -1662 1963 -1610
rect 2499 -2005 3099 -1953
rect 7384 -673 7984 -621
rect 7384 -1021 7984 -969
rect 7383 -1352 7984 -1300
rect 7326 -1599 7378 -1400
rect 7384 -1700 7985 -1648
rect 7142 -1926 7282 -1848
<< metal2 >>
rect 2499 -616 7984 -606
rect 2499 -618 7145 -616
rect 1363 -657 2135 -643
rect 1363 -658 1985 -657
rect 1963 -710 1985 -658
rect 1363 -714 1985 -710
rect 2125 -714 2135 -657
rect 3099 -670 7145 -618
rect 2499 -673 7145 -670
rect 7285 -621 7984 -616
rect 7285 -673 7384 -621
rect 2499 -683 7984 -673
rect 1363 -720 2135 -714
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -897 2355 -887
rect 7133 -969 7984 -959
rect 1363 -1006 2135 -996
rect 1963 -1058 1985 -1006
rect 1363 -1063 1985 -1058
rect 2125 -1063 2135 -1006
rect 7133 -1026 7143 -969
rect 7283 -1021 7384 -969
rect 7283 -1026 7984 -1021
rect 7133 -1036 7984 -1026
rect 1363 -1068 2135 -1063
rect 1363 -1073 2125 -1068
rect 2499 -1164 7293 -1157
rect 2499 -1167 7143 -1164
rect 3099 -1219 7143 -1167
rect 2499 -1221 7143 -1219
rect 7283 -1221 7293 -1164
rect 2499 -1229 7293 -1221
rect 1363 -1257 2355 -1247
rect 1363 -1262 2205 -1257
rect 1963 -1314 2205 -1262
rect 2345 -1314 2355 -1257
rect 1363 -1324 2355 -1314
rect 7133 -1294 7984 -1285
rect 7133 -1351 7143 -1294
rect 7283 -1300 7984 -1294
rect 7283 -1351 7383 -1300
rect 7133 -1352 7383 -1351
rect 7133 -1362 7984 -1352
rect 2499 -1400 7378 -1390
rect 2499 -1405 3177 -1400
rect 1975 -1427 2135 -1417
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 3099 -1457 3177 -1405
rect 3317 -1457 7326 -1400
rect 2499 -1467 7326 -1457
rect 1975 -1494 2135 -1484
rect 1363 -1610 2355 -1600
rect 7326 -1609 7378 -1599
rect 1963 -1662 2205 -1610
rect 1363 -1667 2205 -1662
rect 2345 -1667 2355 -1610
rect 1363 -1672 2355 -1667
rect 7133 -1648 7985 -1638
rect 7133 -1705 7143 -1648
rect 7283 -1700 7384 -1648
rect 7283 -1705 7985 -1700
rect 7133 -1715 7985 -1705
rect 7142 -1848 7282 -1838
rect 7142 -1936 7282 -1926
rect 2499 -1952 3327 -1943
rect 2499 -1953 3177 -1952
rect 3099 -2005 3177 -1953
rect 2499 -2009 3177 -2005
rect 3317 -2009 3327 -1952
rect 2499 -2015 3327 -2009
<< via2 >>
rect 1985 -714 2125 -657
rect 7145 -673 7285 -616
rect 2205 -887 2345 -830
rect 1985 -1063 2125 -1006
rect 7143 -1026 7283 -969
rect 7143 -1221 7283 -1164
rect 2205 -1314 2345 -1257
rect 7143 -1351 7283 -1294
rect 1985 -1484 2125 -1427
rect 3177 -1457 3317 -1400
rect 2205 -1667 2345 -1610
rect 7143 -1705 7283 -1648
rect 7142 -1926 7282 -1848
rect 3177 -2009 3317 -1952
<< metal3 >>
rect 7133 -616 7294 -606
rect 1975 -657 2135 -648
rect 1975 -714 1985 -657
rect 2125 -714 2135 -657
rect 1975 -1006 2135 -714
rect 7133 -673 7145 -616
rect 7285 -673 7294 -616
rect 1975 -1063 1985 -1006
rect 2125 -1063 2135 -1006
rect 1975 -1427 2135 -1063
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 1975 -1494 2135 -1484
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -1257 2355 -887
rect 2195 -1314 2205 -1257
rect 2345 -1314 2355 -1257
rect 2195 -1610 2355 -1314
rect 7133 -969 7294 -673
rect 7133 -1026 7143 -969
rect 7283 -1026 7294 -969
rect 7133 -1164 7294 -1026
rect 7133 -1221 7143 -1164
rect 7283 -1221 7294 -1164
rect 7133 -1294 7294 -1221
rect 7133 -1351 7143 -1294
rect 7283 -1351 7294 -1294
rect 2195 -1667 2205 -1610
rect 2345 -1667 2355 -1610
rect 2195 -1672 2355 -1667
rect 3167 -1400 3327 -1390
rect 3167 -1457 3177 -1400
rect 3317 -1457 3327 -1400
rect 3167 -1952 3327 -1457
rect 7133 -1648 7294 -1351
rect 7133 -1705 7143 -1648
rect 7283 -1705 7294 -1648
rect 7133 -1843 7294 -1705
rect 7132 -1848 7294 -1843
rect 7132 -1926 7142 -1848
rect 7282 -1926 7294 -1848
rect 7132 -1931 7294 -1926
rect 3167 -2009 3177 -1952
rect 3317 -2009 3327 -1952
rect 3167 -2014 3327 -2009
rect 7133 -2015 7294 -1931
use sky130_fd_pr__diode_pw2nd_05v5_37RBXE  sky130_fd_pr__diode_pw2nd_05v5_37RBXE_0
timestamp 1713020003
transform 0 1 7212 -1 0 -1887
box -183 -208 183 208
use sky130_fd_pr__nfet_01v8_MG6U6H  sky130_fd_pr__nfet_01v8_MG6U6H_0
timestamp 1713020003
transform 1 0 7684 0 1 -1500
box -496 -310 496 310
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0
timestamp 1713020003
transform -1 0 2799 0 1 -1705
box -528 -458 528 458
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1
timestamp 1713020003
transform -1 0 2799 0 1 -919
box -528 -458 528 458
use sky130_fd_pr__pfet_01v8_J2L9Q3  sky130_fd_pr__pfet_01v8_J2L9Q3_0
timestamp 1713020003
transform 1 0 7684 0 1 -821
box -496 -319 496 319
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0
timestamp 1713020003
transform 1 0 1663 0 -1 -1462
box -558 -397 558 397
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1
timestamp 1713020003
transform 1 0 1663 0 -1 -858
box -558 -397 558 397
<< labels >>
flabel space 1105 -1255 2221 -461 0 FreeSans 1600 0 0 0 M3
flabel space 2271 -1377 3327 -461 0 FreeSans 1600 0 0 0 M5
flabel space 2271 -2163 3327 -1247 0 FreeSans 1600 0 0 0 M6
flabel metal1 1183 -539 2143 -340 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 1363 -1662 1963 -1610 0 FreeSans 800 0 0 0 out_b
port 2 nsew
flabel metal2 1363 -710 1963 -658 0 FreeSans 800 0 0 0 out
port 3 nsew
flabel space 1105 -1859 2221 -1065 0 FreeSans 1600 0 0 0 M4
flabel metal2 3317 -1467 3773 -1390 0 FreeSans 800 0 0 0 in_b
flabel metal1 2319 -2314 3279 -2115 0 FreeSans 1600 0 0 0 avss
port 4 nsew
flabel space 7224 -538 8184 -340 0 FreeSans 1600 0 0 0 dvdd
port 5 nsew
flabel metal3 7133 -2015 7294 -1926 0 FreeSans 1600 0 0 0 in
port 6 nsew
flabel space 7188 -1810 8180 -1190 0 FreeSans 1600 0 0 0 M1
flabel space 7188 -1140 8180 -502 0 FreeSans 1600 0 0 0 M2
flabel metal1 7040 -2313 8144 -2244 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
<< end >>

magic
tech sky130A
timestamp 1713228232
<< pwell >>
rect -264 -229 264 229
<< mvnmos >>
rect -150 -100 150 100
<< mvndiff >>
rect -179 94 -150 100
rect -179 -94 -173 94
rect -156 -94 -150 94
rect -179 -100 -150 -94
rect 150 94 179 100
rect 150 -94 156 94
rect 173 -94 179 94
rect 150 -100 179 -94
<< mvndiffc >>
rect -173 -94 -156 94
rect 156 -94 173 94
<< mvpsubdiff >>
rect -246 205 246 211
rect -246 188 -192 205
rect 192 188 246 205
rect -246 182 246 188
rect -246 157 -217 182
rect -246 -157 -240 157
rect -223 -157 -217 157
rect 217 157 246 182
rect -246 -182 -217 -157
rect 217 -157 223 157
rect 240 -157 246 157
rect 217 -182 246 -157
rect -246 -188 246 -182
rect -246 -205 -192 -188
rect 192 -205 246 -188
rect -246 -211 246 -205
<< mvpsubdiffcont >>
rect -192 188 192 205
rect -240 -157 -223 157
rect 223 -157 240 157
rect -192 -205 192 -188
<< poly >>
rect -150 136 150 144
rect -150 119 -142 136
rect 142 119 150 136
rect -150 100 150 119
rect -150 -119 150 -100
rect -150 -136 -142 -119
rect 142 -136 150 -119
rect -150 -144 150 -136
<< polycont >>
rect -142 119 142 136
rect -142 -136 142 -119
<< locali >>
rect -240 188 -192 205
rect 192 188 240 205
rect -240 157 -223 188
rect 223 157 240 188
rect -150 119 -142 136
rect 142 119 150 136
rect -173 94 -156 102
rect -173 -102 -156 -94
rect 156 94 173 102
rect 156 -102 173 -94
rect -150 -136 -142 -119
rect 142 -136 150 -119
rect -240 -188 -223 -157
rect 223 -188 240 -157
rect -240 -205 -192 -188
rect 192 -205 240 -188
<< viali >>
rect -142 119 142 136
rect -173 -94 -156 94
rect 156 -94 173 94
rect -142 -136 142 -119
<< metal1 >>
rect -148 136 148 139
rect -148 119 -142 136
rect 142 119 148 136
rect -148 116 148 119
rect -176 94 -153 100
rect -176 -94 -173 94
rect -156 -94 -153 94
rect -176 -100 -153 -94
rect 153 94 176 100
rect 153 -94 156 94
rect 173 -94 176 94
rect 153 -100 176 -94
rect -148 -119 148 -116
rect -148 -136 -142 -119
rect 142 -136 148 -119
rect -148 -139 148 -136
<< properties >>
string FIXED_BBOX -231 -196 231 196
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 2.0 l 3.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

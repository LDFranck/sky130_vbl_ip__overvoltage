magic
tech sky130A
magscale 1 2
timestamp 1712609300
<< nwell >>
rect 19251 1675 19306 1683
rect 17633 1437 19288 1444
rect 19270 1365 19288 1437
<< metal1 >>
rect 17110 2246 19786 2292
rect 17110 1964 17156 2246
rect 17368 1964 17414 2246
rect 17542 1964 17642 2246
rect 19254 1964 19300 2246
rect 19482 1964 19528 2246
rect 19740 1964 19786 2246
rect 17110 1918 19786 1964
rect 17110 1760 17156 1918
rect 17368 1760 17414 1918
rect 17110 1714 17174 1760
rect 17353 1714 17414 1760
rect 17110 1432 17156 1714
rect 17368 1432 17414 1714
rect 17110 1386 17178 1432
rect 17356 1386 17414 1432
rect 17110 1228 17156 1386
rect 17368 1228 17414 1386
rect 5320 1182 16568 1228
rect 5320 900 5366 1182
rect 5578 900 5624 1182
rect 16264 900 16310 1182
rect 16522 900 16568 1182
rect 5320 854 16568 900
rect 5320 696 5366 854
rect 5578 696 5624 854
rect 5320 650 5397 696
rect 5560 650 5624 696
rect 5320 368 5366 650
rect 5578 368 5624 650
rect 5320 322 5393 368
rect 5562 322 5624 368
rect 0 0 200 200
rect 5320 164 5366 322
rect 5578 164 5624 322
rect 5320 118 5394 164
rect 5565 118 5624 164
rect 5320 -164 5366 118
rect 5578 -164 5624 118
rect 0 -400 200 -200
rect 5320 -210 5398 -164
rect 5561 -210 5624 -164
rect 5320 -368 5366 -210
rect 5578 -368 5624 -210
rect 16264 696 16310 854
rect 16522 696 16568 854
rect 16264 650 16339 696
rect 16501 650 16568 696
rect 16264 368 16310 650
rect 16522 368 16568 650
rect 16264 322 16340 368
rect 16504 322 16568 368
rect 16264 164 16310 322
rect 16522 164 16568 322
rect 16264 118 16338 164
rect 16502 118 16568 164
rect 16264 -164 16310 118
rect 16522 -164 16568 118
rect 16264 -210 16343 -164
rect 16499 -210 16568 -164
rect 16264 -368 16310 -210
rect 16522 -368 16568 -210
rect 5320 -414 16568 -368
rect 0 -800 200 -600
rect 5320 -696 5366 -414
rect 5578 -696 5624 -414
rect 16264 -696 16310 -414
rect 16522 -696 16568 -414
rect 5320 -742 16568 -696
rect 17110 1182 17178 1228
rect 17356 1182 17414 1228
rect 17110 900 17156 1182
rect 17368 900 17414 1182
rect 17110 854 17180 900
rect 17356 854 17414 900
rect 17110 696 17156 854
rect 17368 696 17414 854
rect 17110 650 17176 696
rect 17346 650 17414 696
rect 17110 368 17156 650
rect 17368 368 17414 650
rect 17110 322 17178 368
rect 17355 322 17414 368
rect 17110 164 17156 322
rect 17368 164 17414 322
rect 17110 118 17174 164
rect 17353 118 17414 164
rect 17110 -164 17156 118
rect 17368 -164 17414 118
rect 17110 -210 17176 -164
rect 17350 -210 17414 -164
rect 17110 -368 17156 -210
rect 17368 -368 17414 -210
rect 17542 -368 17610 1918
rect 17638 1721 17648 1778
rect 19248 1721 19258 1778
rect 17638 1714 19258 1721
rect 19482 1760 19528 1918
rect 19740 1760 19786 1918
rect 19482 1714 19551 1760
rect 19726 1714 19786 1760
rect 19244 1473 19254 1673
rect 19306 1473 19316 1673
rect 19482 1432 19528 1714
rect 19740 1432 19786 1714
rect 17638 1425 19258 1432
rect 17638 1368 17648 1425
rect 19248 1368 19258 1425
rect 19482 1386 19552 1432
rect 19729 1386 19786 1432
rect 17638 1189 17648 1246
rect 19248 1189 19258 1246
rect 17638 1182 19258 1189
rect 19482 1228 19528 1386
rect 19740 1228 19786 1386
rect 19482 1182 19546 1228
rect 19727 1182 19786 1228
rect 19244 941 19254 1141
rect 19306 941 19316 1141
rect 19482 900 19528 1182
rect 19740 900 19786 1182
rect 17639 893 19259 900
rect 17639 836 17649 893
rect 19249 836 19259 893
rect 19482 854 19549 900
rect 19727 854 19786 900
rect 17638 657 17648 714
rect 19248 657 19258 714
rect 17638 650 19258 657
rect 19482 696 19528 854
rect 19740 696 19786 854
rect 19482 650 19550 696
rect 19726 650 19786 696
rect 19244 409 19254 609
rect 19306 409 19316 609
rect 19482 368 19528 650
rect 19740 368 19786 650
rect 17638 361 19258 368
rect 17638 304 17648 361
rect 19248 304 19258 361
rect 19482 322 19550 368
rect 19728 322 19786 368
rect 17638 125 17648 182
rect 19248 125 19258 182
rect 17638 118 19258 125
rect 19482 164 19528 322
rect 19740 164 19786 322
rect 19482 118 19547 164
rect 19722 118 19786 164
rect 19244 -123 19254 77
rect 19306 -123 19316 77
rect 19482 -164 19528 118
rect 19740 -164 19786 118
rect 17638 -171 19258 -164
rect 17638 -228 17648 -171
rect 19248 -228 19258 -171
rect 19482 -210 19552 -164
rect 19719 -210 19786 -164
rect 19482 -368 19528 -210
rect 19740 -368 19786 -210
rect 17110 -414 19786 -368
rect 17110 -696 17156 -414
rect 17368 -696 17414 -414
rect 17542 -696 17643 -414
rect 19254 -696 19300 -414
rect 19482 -696 19528 -414
rect 19740 -696 19786 -414
rect 17110 -742 19786 -696
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
rect 0 -2400 200 -2200
<< via1 >>
rect 17648 1721 19248 1778
rect 19254 1473 19306 1673
rect 17648 1368 19248 1425
rect 17648 1189 19248 1246
rect 19254 941 19306 1141
rect 17649 836 19249 893
rect 17648 657 19248 714
rect 19254 409 19306 609
rect 17648 304 19248 361
rect 17648 125 19248 182
rect 19254 -123 19306 77
rect 17648 -228 19248 -171
<< metal2 >>
rect 16906 1815 16966 1825
rect 19930 1812 19990 1822
rect 16966 1778 19930 1788
rect 16966 1721 17648 1778
rect 19248 1721 19930 1778
rect 16966 1711 19930 1721
rect 16906 1648 16966 1658
rect 19254 1673 19306 1683
rect 16906 1495 16966 1505
rect 19930 1645 19990 1655
rect 19254 1463 19306 1473
rect 19930 1477 19990 1487
rect 16966 1425 19930 1435
rect 16966 1368 17648 1425
rect 19248 1368 19930 1425
rect 16966 1358 19930 1368
rect 16906 1328 16966 1338
rect 19930 1310 19990 1320
rect 16906 1283 16966 1293
rect 19930 1272 19990 1282
rect 16966 1246 19930 1256
rect 16966 1189 17648 1246
rect 19248 1189 19930 1246
rect 16966 1179 19930 1189
rect 16906 1116 16966 1126
rect 19254 1141 19306 1151
rect 16906 957 16966 967
rect 19930 1105 19990 1115
rect 19254 931 19306 941
rect 19930 948 19990 958
rect 16966 893 19930 903
rect 16966 836 17649 893
rect 19249 836 19930 893
rect 16966 826 19930 836
rect 16906 790 16966 800
rect 19930 781 19990 791
rect 16906 752 16966 762
rect 19930 741 19990 751
rect 16966 714 19930 724
rect 16966 657 17648 714
rect 19248 657 19930 714
rect 16966 647 19930 657
rect 16906 585 16966 595
rect 19254 609 19306 619
rect 16906 429 16966 439
rect 19930 574 19990 584
rect 19254 399 19306 409
rect 19930 424 19990 434
rect 16966 361 19930 371
rect 16966 304 17648 361
rect 19248 304 19930 361
rect 16966 294 19930 304
rect 16906 262 16966 272
rect 19930 257 19990 267
rect 16906 222 16966 232
rect 19930 216 19990 226
rect 16966 182 19930 192
rect 16966 125 17648 182
rect 19248 125 19930 182
rect 16966 115 19930 125
rect 16906 55 16966 65
rect 19254 77 19306 87
rect 16906 -111 16966 -101
rect 19930 49 19990 59
rect 19254 -133 19306 -123
rect 19930 -116 19990 -106
rect 16966 -171 19930 -161
rect 16966 -228 17648 -171
rect 19248 -228 19930 -171
rect 16966 -238 19930 -228
rect 16906 -278 16966 -268
rect 19930 -283 19990 -273
<< via2 >>
rect 16906 1658 16966 1815
rect 16906 1338 16966 1495
rect 19930 1655 19990 1812
rect 19930 1320 19990 1477
rect 16906 1126 16966 1283
rect 16906 800 16966 957
rect 19930 1115 19990 1272
rect 19930 791 19990 948
rect 16906 595 16966 752
rect 16906 272 16966 429
rect 19930 584 19990 741
rect 19930 267 19990 424
rect 16906 65 16966 222
rect 16906 -268 16966 -111
rect 19930 59 19990 216
rect 19930 -273 19990 -116
<< metal3 >>
rect 16896 1815 16976 1836
rect 16896 1658 16906 1815
rect 16966 1658 16976 1815
rect 16896 1495 16976 1658
rect 16896 1338 16906 1495
rect 16966 1338 16976 1495
rect 16896 1283 16976 1338
rect 16896 1126 16906 1283
rect 16966 1126 16976 1283
rect 16896 957 16976 1126
rect 16896 800 16906 957
rect 16966 800 16976 957
rect 16896 752 16976 800
rect 16896 595 16906 752
rect 16966 595 16976 752
rect 16896 429 16976 595
rect 16896 272 16906 429
rect 16966 272 16976 429
rect 16896 222 16976 272
rect 16896 65 16906 222
rect 16966 65 16976 222
rect 16896 -111 16976 65
rect 16896 -268 16906 -111
rect 16966 -268 16976 -111
rect 16896 -742 16976 -268
rect 19920 1812 20000 1833
rect 19920 1655 19930 1812
rect 19990 1655 20000 1812
rect 19920 1477 20000 1655
rect 19920 1320 19930 1477
rect 19990 1320 20000 1477
rect 19920 1272 20000 1320
rect 19920 1115 19930 1272
rect 19990 1115 20000 1272
rect 19920 948 20000 1115
rect 19920 791 19930 948
rect 19990 791 20000 948
rect 19920 741 20000 791
rect 19920 584 19930 741
rect 19990 584 20000 741
rect 19920 424 20000 584
rect 19920 267 19930 424
rect 19990 267 20000 424
rect 19920 216 20000 267
rect 19920 59 19930 216
rect 19990 59 20000 216
rect 19920 -116 20000 59
rect 19920 -273 19930 -116
rect 19990 -273 20000 -116
rect 19920 -742 20000 -273
rect 20060 -744 20140 1833
use trans_gate  x1
timestamp 1712344797
transform 1 0 3352 0 1 -2005
box 0 -2052 3413 715
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[0]
timestamp 1712597941
transform 1 0 15047 0 1 -2072
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[1]
timestamp 1712597941
transform 1 0 15047 0 1 -3364
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[0]
timestamp 1712597941
transform 1 0 15047 0 1 -2718
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[1]
timestamp 1712597941
transform 1 0 15047 0 1 -4010
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[0]
timestamp 1712343889
transform 1 0 18448 0 1 1041
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[1]
timestamp 1712343889
transform 1 0 18448 0 1 509
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM4[0]
timestamp 1712343889
transform 1 0 10944 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM4[1]
timestamp 1712343889
transform 1 0 10944 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[0]
timestamp 1712343889
transform 1 0 18448 0 1 1573
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[1]
timestamp 1712343889
transform 1 0 18448 0 1 -23
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[0]
timestamp 1712343889
transform 1 0 7458 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[1]
timestamp 1712343889
transform 1 0 7458 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[2]
timestamp 1712343889
transform 1 0 14430 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[3]
timestamp 1712343889
transform 1 0 14430 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1712343889
transform 1 0 17953 0 1 -1841
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_697RXD  XM8
timestamp 1712343889
transform 1 0 17953 0 1 -2906
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1712343889
transform 1 0 19502 0 1 -1649
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1712343889
transform 1 0 19402 0 1 -3126
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1712343889
transform 1 0 10757 0 1 -2114
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1712343889
transform 1 0 10738 0 1 -1380
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1712343889
transform 1 0 12457 0 1 -2895
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1712343889
transform 1 0 12449 0 1 -3612
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1712343889
transform 1 0 16006 0 1 2117
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1712343889
transform 1 0 14718 0 1 2136
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1712343889
transform 1 0 17483 0 1 -3659
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1712343889
transform 1 0 7558 0 1 -1447
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1712343889
transform 1 0 7558 0 1 -2201
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[0]
timestamp 1712344493
transform 1 0 17262 0 1 2105
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[1]
timestamp 1712344493
transform 1 0 17262 0 1 1573
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[2]
timestamp 1712344493
transform 1 0 17262 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[3]
timestamp 1712344493
transform 1 0 17262 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712344493
transform 1 0 17262 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712344493
transform 1 0 17262 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712344493
transform 1 0 19634 0 1 2105
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712344493
transform 1 0 19634 0 1 1573
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712344493
transform 1 0 19634 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712344493
transform 1 0 19634 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712344493
transform 1 0 19634 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712344493
transform 1 0 19634 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712344493
transform 1 0 5472 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712344493
transform 1 0 5472 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712344493
transform 1 0 5472 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712344493
transform 1 0 5472 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[16]
timestamp 1712344493
transform 1 0 16416 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[17]
timestamp 1712344493
transform 1 0 16416 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[18]
timestamp 1712344493
transform 1 0 16416 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[19]
timestamp 1712344493
transform 1 0 16416 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[0]
timestamp 1712343889
transform 1 0 18448 0 1 2105
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[1]
timestamp 1712343889
transform 1 0 18448 0 1 -555
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712344493
transform 1 0 7458 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712344493
transform 1 0 10944 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712344493
transform 1 0 14430 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712344493
transform 1 0 7458 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712344493
transform 1 0 10944 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712344493
transform 1 0 14430 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712600458
transform 1 0 13709 0 1 -1456
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712600458
transform 1 0 13709 0 1 -4626
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712600458
transform 1 0 16385 0 1 -1456
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712600458
transform 1 0 16385 0 1 -4626
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712599722
transform 1 0 15047 0 1 -1456
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712599722
transform 1 0 15047 0 1 -4626
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712597941
transform 1 0 13709 0 1 -2072
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712597941
transform 1 0 13709 0 1 -2718
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712597941
transform 1 0 13709 0 1 -3364
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712597941
transform 1 0 13709 0 1 -4010
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[4]
timestamp 1712597941
transform 1 0 16385 0 1 -2072
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[5]
timestamp 1712597941
transform 1 0 16385 0 1 -2718
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[6]
timestamp 1712597941
transform 1 0 16385 0 1 -3364
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[7]
timestamp 1712597941
transform 1 0 16385 0 1 -4010
box -328 -388 328 388
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 dvdd
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 out
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 vref
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 vin
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 ena
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 ibias
port 5 nsew
flabel metal1 0 -2400 200 -2200 0 FreeSans 256 0 0 0 vss
port 6 nsew
<< end >>

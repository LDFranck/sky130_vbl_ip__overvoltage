magic
tech sky130A
timestamp 1711994542
<< pwell >>
rect -498 -155 498 155
<< nmos >>
rect -400 -50 400 50
<< ndiff >>
rect -429 44 -400 50
rect -429 -44 -423 44
rect -406 -44 -400 44
rect -429 -50 -400 -44
rect 400 44 429 50
rect 400 -44 406 44
rect 423 -44 429 44
rect 400 -50 429 -44
<< ndiffc >>
rect -423 -44 -406 44
rect 406 -44 423 44
<< psubdiff >>
rect -480 120 -432 137
rect 432 120 480 137
rect -480 89 -463 120
rect 463 89 480 120
rect -480 -120 -463 -89
rect 463 -120 480 -89
rect -480 -137 -432 -120
rect 432 -137 480 -120
<< psubdiffcont >>
rect -432 120 432 137
rect -480 -89 -463 89
rect 463 -89 480 89
rect -432 -137 432 -120
<< poly >>
rect -400 86 400 94
rect -400 69 -392 86
rect 392 69 400 86
rect -400 50 400 69
rect -400 -69 400 -50
rect -400 -86 -392 -69
rect 392 -86 400 -69
rect -400 -94 400 -86
<< polycont >>
rect -392 69 392 86
rect -392 -86 392 -69
<< locali >>
rect -480 120 -432 137
rect 432 120 480 137
rect -480 89 -463 120
rect 463 89 480 120
rect -400 69 -392 86
rect 392 69 400 86
rect -423 44 -406 52
rect -423 -52 -406 -44
rect 406 44 423 52
rect 406 -52 423 -44
rect -400 -86 -392 -69
rect 392 -86 400 -69
rect -480 -120 -463 -89
rect 463 -120 480 -89
rect -480 -137 -432 -120
rect 432 -137 480 -120
<< viali >>
rect -392 69 392 86
rect -423 -44 -406 44
rect 406 -44 423 44
rect -392 -86 392 -69
<< metal1 >>
rect -398 86 398 89
rect -398 69 -392 86
rect 392 69 398 86
rect -398 66 398 69
rect -426 44 -403 50
rect -426 -44 -423 44
rect -406 -44 -403 44
rect -426 -50 -403 -44
rect 403 44 426 50
rect 403 -44 406 44
rect 423 -44 426 44
rect 403 -50 426 -44
rect -398 -69 398 -66
rect -398 -86 -392 -69
rect 392 -86 398 -69
rect -398 -89 398 -86
<< properties >>
string FIXED_BBOX -471 -128 471 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 8.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

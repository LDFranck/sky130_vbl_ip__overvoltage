magic
tech sky130A
magscale 1 2
timestamp 1713221383
<< metal1 >>
rect -3578 12199 -3568 12373
rect -3448 12199 -3438 12373
rect -3568 9295 -3448 12199
rect -3388 10589 -3378 10763
rect -3258 10589 -3248 10763
rect -3578 8993 -3568 9295
rect -3448 8993 -3438 9295
rect -3378 8539 -3258 10589
rect -3198 8979 -3188 9153
rect -3068 8979 -3058 9153
rect -3388 8237 -3378 8539
rect -3258 8237 -3248 8539
rect -3188 6649 -3068 8979
rect -3008 7369 -2998 7543
rect -2878 7369 -2868 7543
rect -3198 6347 -3188 6649
rect -3068 6347 -3058 6649
rect -2998 5893 -2878 7369
rect -3008 5591 -2998 5893
rect -2878 5591 -2868 5893
rect -2818 5759 -2808 5933
rect -2688 5759 -2678 5933
rect -2808 4381 -2688 5759
rect -2818 4079 -2808 4381
rect -2688 4079 -2678 4381
rect -2628 4149 -2618 4323
rect -2498 4149 -2488 4323
rect -2618 4003 -2498 4149
rect -2628 3701 -2618 4003
rect -2498 3701 -2488 4003
rect -3578 2189 -3568 2491
rect -3448 2189 -3438 2491
rect -3568 1157 -3448 2189
rect -3578 983 -3568 1157
rect -3448 983 -3438 1157
<< via1 >>
rect -3568 12199 -3448 12373
rect -3378 10589 -3258 10763
rect -3568 8993 -3448 9295
rect -3188 8979 -3068 9153
rect -3378 8237 -3258 8539
rect -2998 7369 -2878 7543
rect -3188 6347 -3068 6649
rect -2998 5591 -2878 5893
rect -2808 5759 -2688 5933
rect -2808 4079 -2688 4381
rect -2618 4149 -2498 4323
rect -2618 3701 -2498 4003
rect -3568 2189 -3448 2491
rect -3568 983 -3448 1157
<< metal2 >>
rect -3568 12373 -3448 12383
rect -3448 12253 -2619 12373
rect -3568 12189 -3448 12199
rect -3378 10763 -3258 10773
rect -3258 10643 -2619 10763
rect -3378 10579 -3258 10589
rect -3568 9295 -3448 9305
rect -3568 8983 -3448 8993
rect -3188 9153 -3068 9163
rect -3068 9033 -2619 9153
rect -3188 8969 -3068 8979
rect -3378 8539 -3258 8549
rect -3448 8237 -3378 8539
rect -3378 8227 -3258 8237
rect -3568 7783 -3448 7793
rect -3568 7471 -3448 7481
rect -2998 7543 -2878 7553
rect -2878 7423 -2619 7543
rect -2998 7359 -2878 7369
rect -3378 7027 -3258 7037
rect -3448 6725 -3378 7027
rect -3378 6715 -3258 6725
rect -3188 6649 -3068 6659
rect -3448 6347 -3188 6649
rect -3188 6337 -3068 6347
rect -2808 5933 -2688 5943
rect -2998 5893 -2878 5903
rect -3448 5591 -2998 5893
rect -2688 5813 -2619 5933
rect -2808 5749 -2688 5759
rect -2998 5581 -2878 5591
rect -3188 5515 -3068 5525
rect -3448 5213 -3188 5515
rect -3188 5203 -3068 5213
rect -2998 4759 -2878 4769
rect -3448 4457 -2998 4759
rect -2998 4447 -2878 4457
rect -2808 4381 -2688 4391
rect -3448 4079 -2808 4381
rect -2618 4323 -2498 4333
rect -2618 4139 -2498 4149
rect -2808 4069 -2688 4079
rect -2618 4003 -2498 4013
rect -3448 3701 -2618 4003
rect -2618 3691 -2498 3701
rect -2808 3625 -2688 3635
rect -3448 3323 -2808 3625
rect -2808 3313 -2688 3323
rect -2618 3247 -2498 3257
rect -3448 2945 -2618 3247
rect -2618 2935 -2498 2945
rect -3448 2593 -2619 2713
rect -3568 2491 -3448 2501
rect -3568 2179 -3448 2189
rect -3378 2113 -3258 2123
rect -3448 1811 -3378 2113
rect -3378 1801 -3258 1811
rect -3568 1735 -3448 1745
rect -3568 1423 -3448 1433
rect -3568 1157 -3448 1167
rect -3448 983 -2619 1103
rect -3568 973 -3448 983
<< via2 >>
rect -3568 7481 -3448 7783
rect -3378 6725 -3258 7027
rect -3188 5213 -3068 5515
rect -2998 4457 -2878 4759
rect -2808 3323 -2688 3625
rect -2618 2945 -2498 3247
rect -3378 1811 -3258 2113
rect -3568 1433 -3448 1735
<< metal3 >>
rect -3578 12199 -3568 12373
rect -3448 12199 -3438 12373
rect -3568 7788 -3448 12199
rect -3388 10589 -3378 10763
rect -3258 10589 -3248 10763
rect -3578 7783 -3438 7788
rect -3578 7481 -3568 7783
rect -3448 7481 -3438 7783
rect -3578 7476 -3438 7481
rect -3378 7032 -3258 10589
rect -3198 8979 -3188 9153
rect -3068 8979 -3058 9153
rect -3388 7027 -3248 7032
rect -3388 6725 -3378 7027
rect -3258 6725 -3248 7027
rect -3388 6720 -3248 6725
rect -3188 5520 -3068 8979
rect -3008 7369 -2998 7543
rect -2878 7369 -2868 7543
rect -3198 5515 -3058 5520
rect -3198 5213 -3188 5515
rect -3068 5213 -3058 5515
rect -3198 5208 -3058 5213
rect -2998 4764 -2878 7369
rect -2818 5759 -2808 5933
rect -2688 5759 -2678 5933
rect -3008 4759 -2868 4764
rect -3008 4457 -2998 4759
rect -2878 4457 -2868 4759
rect -3008 4452 -2868 4457
rect -2808 3630 -2688 5759
rect -2628 4149 -2618 4323
rect -2498 4149 -2488 4323
rect -2818 3625 -2678 3630
rect -2818 3323 -2808 3625
rect -2688 3323 -2678 3625
rect -2818 3318 -2678 3323
rect -2618 3252 -2498 4149
rect -2628 3247 -2488 3252
rect -2628 2945 -2618 3247
rect -2498 2945 -2488 3247
rect -2628 2940 -2488 2945
rect -3388 2539 -3378 2713
rect -3258 2539 -3248 2713
rect -3378 2118 -3258 2539
rect -3388 2113 -3248 2118
rect -3388 1811 -3378 2113
rect -3258 1811 -3248 2113
rect -3388 1806 -3248 1811
rect -3578 1735 -3438 1740
rect -3578 1433 -3568 1735
rect -3448 1433 -3438 1735
rect -3578 1428 -3438 1433
rect -3568 1157 -3448 1428
rect -3578 983 -3568 1157
rect -3448 983 -3438 1157
<< via3 >>
rect -3568 12199 -3448 12373
rect -3378 10589 -3258 10763
rect -3188 8979 -3068 9153
rect -2998 7369 -2878 7543
rect -2808 5759 -2688 5933
rect -2618 4149 -2498 4323
rect -3378 2539 -3258 2713
rect -3568 983 -3448 1157
<< metal4 >>
rect -3569 12373 -3447 12374
rect -3569 12199 -3568 12373
rect -3448 12364 -3447 12373
rect -3448 12262 -2519 12364
rect -3448 12199 -3447 12262
rect -3569 12198 -3447 12199
rect -3379 10763 -3257 10764
rect -3379 10589 -3378 10763
rect -3258 10754 -3257 10763
rect -3258 10652 -2519 10754
rect -3258 10589 -3257 10652
rect -3379 10588 -3257 10589
rect -3189 9153 -3067 9154
rect -3189 8979 -3188 9153
rect -3068 9144 -3067 9153
rect -3068 9042 -2519 9144
rect -3068 8979 -3067 9042
rect -3189 8978 -3067 8979
rect -2999 7543 -2877 7544
rect -2999 7369 -2998 7543
rect -2878 7534 -2877 7543
rect -2878 7432 -2519 7534
rect -2878 7369 -2877 7432
rect -2999 7368 -2877 7369
rect -2809 5933 -2687 5934
rect -2809 5759 -2808 5933
rect -2688 5924 -2687 5933
rect -2688 5822 -2519 5924
rect -2688 5759 -2687 5822
rect -2809 5758 -2687 5759
rect -2619 4323 -2497 4324
rect -2619 4149 -2618 4323
rect -2498 4149 -2497 4323
rect -2619 4148 -2497 4149
rect -3379 2713 -3257 2714
rect -3379 2539 -3378 2713
rect -3258 2704 -3257 2713
rect -3258 2602 -2519 2704
rect -3258 2539 -3257 2602
rect -3379 2538 -3257 2539
rect -3569 1157 -3447 1158
rect -3569 983 -3568 1157
rect -3448 1094 -3447 1157
rect -3448 992 -2519 1094
rect -3448 983 -3447 992
rect -3569 982 -3447 983
<< end >>

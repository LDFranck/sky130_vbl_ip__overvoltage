magic
tech sky130A
timestamp 1712599722
<< pwell >>
rect -564 -179 564 179
<< mvnmos >>
rect -450 -50 450 50
<< mvndiff >>
rect -479 44 -450 50
rect -479 -44 -473 44
rect -456 -44 -450 44
rect -479 -50 -450 -44
rect 450 44 479 50
rect 450 -44 456 44
rect 473 -44 479 44
rect 450 -50 479 -44
<< mvndiffc >>
rect -473 -44 -456 44
rect 456 -44 473 44
<< mvpsubdiff >>
rect -546 155 546 161
rect -546 138 -492 155
rect 492 138 546 155
rect -546 132 546 138
rect -546 107 -517 132
rect -546 -107 -540 107
rect -523 -107 -517 107
rect 517 107 546 132
rect -546 -132 -517 -107
rect 517 -107 523 107
rect 540 -107 546 107
rect 517 -132 546 -107
rect -546 -138 546 -132
rect -546 -155 -492 -138
rect 492 -155 546 -138
rect -546 -161 546 -155
<< mvpsubdiffcont >>
rect -492 138 492 155
rect -540 -107 -523 107
rect 523 -107 540 107
rect -492 -155 492 -138
<< poly >>
rect -450 86 450 94
rect -450 69 -442 86
rect 442 69 450 86
rect -450 50 450 69
rect -450 -69 450 -50
rect -450 -86 -442 -69
rect 442 -86 450 -69
rect -450 -94 450 -86
<< polycont >>
rect -442 69 442 86
rect -442 -86 442 -69
<< locali >>
rect -540 138 -492 155
rect 492 138 540 155
rect -540 107 -523 138
rect 523 107 540 138
rect -450 69 -442 86
rect 442 69 450 86
rect -473 44 -456 52
rect -473 -52 -456 -44
rect 456 44 473 52
rect 456 -52 473 -44
rect -450 -86 -442 -69
rect 442 -86 450 -69
rect -540 -138 -523 -107
rect 523 -138 540 -107
rect -540 -155 -492 -138
rect 492 -155 540 -138
<< viali >>
rect -442 69 442 86
rect -473 -44 -456 44
rect 456 -44 473 44
rect -442 -86 442 -69
<< metal1 >>
rect -448 86 448 89
rect -448 69 -442 86
rect 442 69 448 86
rect -448 66 448 69
rect -476 44 -453 50
rect -476 -44 -473 44
rect -456 -44 -453 44
rect -476 -50 -453 -44
rect 453 44 476 50
rect 453 -44 456 44
rect 473 -44 476 44
rect 453 -50 476 -44
rect -448 -69 448 -66
rect -448 -86 -442 -69
rect 442 -86 448 -69
rect -448 -89 448 -86
<< properties >>
string FIXED_BBOX -531 -146 531 146
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 9 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

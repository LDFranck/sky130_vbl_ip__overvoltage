magic
tech sky130A
timestamp 1712150472
<< pwell >>
rect -498 -170 498 170
<< nmos >>
rect -400 -65 400 65
<< ndiff >>
rect -429 59 -400 65
rect -429 -59 -423 59
rect -406 -59 -400 59
rect -429 -65 -400 -59
rect 400 59 429 65
rect 400 -59 406 59
rect 423 -59 429 59
rect 400 -65 429 -59
<< ndiffc >>
rect -423 -59 -406 59
rect 406 -59 423 59
<< psubdiff >>
rect -480 135 -432 152
rect 432 135 480 152
rect -480 104 -463 135
rect 463 104 480 135
rect -480 -135 -463 -104
rect 463 -135 480 -104
rect -480 -152 -432 -135
rect 432 -152 480 -135
<< psubdiffcont >>
rect -432 135 432 152
rect -480 -104 -463 104
rect 463 -104 480 104
rect -432 -152 432 -135
<< poly >>
rect -400 101 400 109
rect -400 84 -392 101
rect 392 84 400 101
rect -400 65 400 84
rect -400 -84 400 -65
rect -400 -101 -392 -84
rect 392 -101 400 -84
rect -400 -109 400 -101
<< polycont >>
rect -392 84 392 101
rect -392 -101 392 -84
<< locali >>
rect -480 135 -432 152
rect 432 135 480 152
rect -480 104 -463 135
rect 463 104 480 135
rect -400 84 -392 101
rect 392 84 400 101
rect -423 59 -406 67
rect -423 -67 -406 -59
rect 406 59 423 67
rect 406 -67 423 -59
rect -400 -101 -392 -84
rect 392 -101 400 -84
rect -480 -135 -463 -104
rect 463 -135 480 -104
rect -480 -152 -432 -135
rect 432 -152 480 -135
<< viali >>
rect -392 84 392 101
rect -423 -59 -406 59
rect 406 -59 423 59
rect -392 -101 392 -84
<< metal1 >>
rect -398 101 398 104
rect -398 84 -392 101
rect 392 84 398 101
rect -398 81 398 84
rect -426 59 -403 65
rect -426 -59 -423 59
rect -406 -59 -403 59
rect -426 -65 -403 -59
rect 403 59 426 65
rect 403 -59 406 59
rect 423 -59 426 59
rect 403 -65 426 -59
rect -398 -84 398 -81
rect -398 -101 -392 -84
rect 392 -101 398 -84
rect -398 -104 398 -101
<< properties >>
string FIXED_BBOX -471 -143 471 143
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.3 l 8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713118140
<< nwell >>
rect -18431 17037 7811 17047
rect -18431 16761 7813 17037
rect -18431 -3615 -18145 16761
rect 7525 8905 7813 16761
rect 7525 8619 10386 8905
rect 7622 8610 10386 8619
rect 10100 -3615 10386 8610
rect -18431 -3901 10386 -3615
use comp_hyst  comp_hyst_0
timestamp 1713115829
transform 1 0 8609 0 1 10759
box 1667 -5363 16947 2564
use level_shifter  level_shifter_0
timestamp 1713117387
transform 1 0 6519 0 1 8816
box 1105 -2314 8184 -340
use level_shifter  level_shifter_1
timestamp 1713117387
transform 1 0 6519 0 1 6624
box 1105 -2314 8184 -340
use level_shifter  level_shifter_2
timestamp 1713117387
transform 1 0 6529 0 1 4422
box 1105 -2314 8184 -340
use level_shifter  level_shifter_3
timestamp 1713117387
transform 1 0 6551 0 1 2240
box 1105 -2314 8184 -340
use multiplexer  multiplexer_0
timestamp 1713115829
transform 1 0 -1139 0 1 -203
box -199 -135 8108 13095
use voltage_divider  voltage_divider_0
timestamp 1713115829
transform 1 0 -16349 0 1 -2158
box -1259 -1438 14153 19128
<< end >>

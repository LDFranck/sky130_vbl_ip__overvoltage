magic
tech sky130A
magscale 1 2
timestamp 1712672837
<< nwell >>
rect 15899 1675 15954 1683
rect 14281 1437 15936 1444
rect 15918 1365 15936 1437
<< metal1 >>
rect 13758 2246 16434 2292
rect 13758 1964 13804 2246
rect 14016 1964 14062 2246
rect 14190 1964 14290 2246
rect 15902 1964 15948 2246
rect 16130 1964 16176 2246
rect 16388 1964 16434 2246
rect 13758 1918 16434 1964
rect 13758 1760 13804 1918
rect 14016 1760 14062 1918
rect 13758 1714 13822 1760
rect 14001 1714 14062 1760
rect 13758 1432 13804 1714
rect 14016 1432 14062 1714
rect 13758 1386 13826 1432
rect 14004 1386 14062 1432
rect 13758 1228 13804 1386
rect 14016 1228 14062 1386
rect 1811 1182 13059 1228
rect 1811 900 1857 1182
rect 2069 900 2115 1182
rect 2265 900 2343 1182
rect 5555 900 5601 1182
rect 5751 900 5829 1182
rect 9041 900 9087 1182
rect 9237 900 9315 1182
rect 12527 900 12573 1182
rect 12755 900 12801 1182
rect 13013 900 13059 1182
rect 1811 854 13059 900
rect 1811 696 1857 854
rect 2069 696 2115 854
rect 1811 650 1888 696
rect 2051 650 2115 696
rect 1811 368 1857 650
rect 2069 368 2115 650
rect 1811 322 1884 368
rect 2053 322 2115 368
rect 1811 164 1857 322
rect 2069 164 2115 322
rect 1811 118 1885 164
rect 2056 118 2115 164
rect 1811 -164 1857 118
rect 2069 -164 2115 118
rect 1811 -210 1889 -164
rect 2052 -210 2115 -164
rect 1811 -368 1857 -210
rect 2069 -368 2115 -210
rect 2265 -368 2311 854
rect 2339 657 2349 713
rect 5549 657 5559 713
rect 2339 650 5559 657
rect 5545 409 5555 609
rect 5607 409 5617 609
rect 2339 361 5559 368
rect 2339 305 2349 361
rect 5549 305 5559 361
rect 2339 125 2349 181
rect 5549 125 5559 181
rect 2339 118 5559 125
rect 5545 -123 5555 77
rect 5607 -123 5617 77
rect 2339 -171 5559 -164
rect 2339 -227 2349 -171
rect 5549 -227 5559 -171
rect 5751 -368 5797 854
rect 5825 657 5835 713
rect 9035 657 9087 713
rect 5825 650 9087 657
rect 9041 609 9087 650
rect 9041 368 9087 409
rect 5825 361 9087 368
rect 5825 305 5835 361
rect 9035 305 9087 361
rect 5825 125 5835 181
rect 9035 125 9087 181
rect 5825 118 9087 125
rect 9041 77 9087 118
rect 9041 -164 9087 -123
rect 5825 -171 9087 -164
rect 5825 -227 5835 -171
rect 9035 -227 9087 -171
rect 9237 -368 9283 854
rect 9311 657 9321 713
rect 12521 657 12531 713
rect 9311 650 12531 657
rect 12755 696 12801 854
rect 13013 696 13059 854
rect 12755 650 12830 696
rect 12992 650 13059 696
rect 12517 409 12527 609
rect 12579 409 12589 609
rect 12755 368 12801 650
rect 13013 368 13059 650
rect 9311 361 12531 368
rect 9311 305 9321 361
rect 12521 305 12531 361
rect 12755 322 12831 368
rect 12995 322 13059 368
rect 9311 125 9321 181
rect 12521 125 12531 181
rect 9311 118 12531 125
rect 12755 164 12801 322
rect 13013 164 13059 322
rect 12755 118 12829 164
rect 12993 118 13059 164
rect 12517 -123 12527 77
rect 12579 -123 12589 77
rect 12755 -164 12801 118
rect 13013 -164 13059 118
rect 9311 -171 12531 -164
rect 9311 -227 9321 -171
rect 12521 -227 12531 -171
rect 12755 -210 12834 -164
rect 12990 -210 13059 -164
rect 12755 -368 12801 -210
rect 13013 -368 13059 -210
rect 1811 -414 13059 -368
rect 1811 -696 1857 -414
rect 2069 -696 2115 -414
rect 2265 -696 2343 -414
rect 5555 -696 5601 -414
rect 5751 -696 5829 -414
rect 9041 -696 9087 -414
rect 9237 -696 9315 -414
rect 12527 -696 12573 -414
rect 12755 -696 12801 -414
rect 13013 -696 13059 -414
rect 1811 -742 13059 -696
rect 13758 1182 13826 1228
rect 14004 1182 14062 1228
rect 13758 900 13804 1182
rect 14016 900 14062 1182
rect 13758 854 13828 900
rect 14004 854 14062 900
rect 13758 696 13804 854
rect 14016 696 14062 854
rect 13758 650 13824 696
rect 13994 650 14062 696
rect 13758 368 13804 650
rect 14016 368 14062 650
rect 13758 322 13826 368
rect 14003 322 14062 368
rect 13758 164 13804 322
rect 14016 164 14062 322
rect 13758 118 13822 164
rect 14001 118 14062 164
rect 13758 -164 13804 118
rect 14016 -164 14062 118
rect 13758 -210 13824 -164
rect 13998 -210 14062 -164
rect 13758 -368 13804 -210
rect 14016 -368 14062 -210
rect 14190 -368 14258 1918
rect 14286 1721 14296 1778
rect 15896 1721 15906 1778
rect 14286 1714 15906 1721
rect 16130 1760 16176 1918
rect 16388 1760 16434 1918
rect 16130 1714 16199 1760
rect 16374 1714 16434 1760
rect 15892 1473 15902 1673
rect 15954 1473 15964 1673
rect 16130 1432 16176 1714
rect 16388 1432 16434 1714
rect 14286 1425 15906 1432
rect 14286 1368 14296 1425
rect 15896 1368 15906 1425
rect 16130 1386 16200 1432
rect 16377 1386 16434 1432
rect 14286 1189 14296 1246
rect 15896 1189 15948 1246
rect 14286 1182 15948 1189
rect 15902 1140 15948 1182
rect 16130 1228 16176 1386
rect 16388 1228 16434 1386
rect 16130 1182 16194 1228
rect 16375 1182 16434 1228
rect 15902 900 15948 941
rect 14287 893 15948 900
rect 14287 836 14297 893
rect 15897 836 15948 893
rect 16130 900 16176 1182
rect 16388 900 16434 1182
rect 16130 854 16197 900
rect 16375 854 16434 900
rect 14286 657 14296 714
rect 15896 657 15948 714
rect 14286 650 15948 657
rect 15902 609 15948 650
rect 16130 696 16176 854
rect 16388 696 16434 854
rect 16130 650 16198 696
rect 16374 650 16434 696
rect 15902 368 15948 409
rect 14286 361 15948 368
rect 14286 304 14296 361
rect 15896 304 15948 361
rect 16130 368 16176 650
rect 16388 368 16434 650
rect 16130 322 16198 368
rect 16376 322 16434 368
rect 14286 125 14296 182
rect 15896 125 15906 182
rect 14286 118 15906 125
rect 16130 164 16176 322
rect 16388 164 16434 322
rect 16130 118 16195 164
rect 16370 118 16434 164
rect 15892 -123 15902 77
rect 15954 -123 15964 77
rect 16130 -164 16176 118
rect 16388 -164 16434 118
rect 14286 -171 15906 -164
rect 14286 -228 14296 -171
rect 15896 -228 15906 -171
rect 16130 -210 16200 -164
rect 16367 -210 16434 -164
rect 16130 -368 16176 -210
rect 16388 -368 16434 -210
rect 20126 -329 20326 -129
rect 13758 -414 16434 -368
rect 13758 -696 13804 -414
rect 14016 -696 14062 -414
rect 14190 -696 14291 -414
rect 15902 -696 15948 -414
rect 16130 -696 16176 -414
rect 16388 -696 16434 -414
rect 13758 -742 16434 -696
rect 20126 -729 20326 -529
rect 20126 -1129 20326 -929
rect 20126 -1529 20326 -1329
rect 20126 -1929 20326 -1729
rect 20126 -2329 20326 -2129
rect 20126 -2729 20326 -2529
<< via1 >>
rect 2349 657 5549 713
rect 5555 409 5607 609
rect 2349 305 5549 361
rect 2349 125 5549 181
rect 5555 -123 5607 77
rect 2349 -227 5549 -171
rect 5835 657 9035 713
rect 5835 305 9035 361
rect 5835 125 9035 181
rect 5835 -227 9035 -171
rect 9321 657 12521 713
rect 12527 409 12579 609
rect 9321 305 12521 361
rect 9321 125 12521 181
rect 12527 -123 12579 77
rect 9321 -227 12521 -171
rect 14296 1721 15896 1778
rect 15902 1473 15954 1673
rect 14296 1368 15896 1425
rect 14296 1189 15896 1246
rect 14297 836 15897 893
rect 14296 657 15896 714
rect 14296 304 15896 361
rect 14296 125 15896 182
rect 15902 -123 15954 77
rect 14296 -228 15896 -171
<< metal2 >>
rect 13457 1781 16735 1791
rect 13614 1778 16578 1781
rect 13614 1721 14296 1778
rect 15896 1721 16578 1778
rect 13457 1711 16735 1721
rect 15902 1673 16974 1683
rect 15954 1473 16823 1673
rect 16964 1473 16974 1673
rect 15902 1463 16974 1473
rect 13457 1425 16735 1435
rect 13614 1368 14296 1425
rect 15896 1368 16578 1425
rect 13614 1365 16578 1368
rect 13457 1355 16735 1365
rect 13457 1249 16735 1259
rect 13614 1246 16578 1249
rect 13614 1189 14296 1246
rect 15896 1189 16578 1246
rect 13457 1179 16735 1189
rect 13457 893 16735 903
rect 5504 833 13457 836
rect 13614 836 14297 893
rect 15897 836 16578 893
rect 13614 833 16578 836
rect 5504 826 16735 833
rect 5661 766 12471 826
rect 12628 823 16735 826
rect 12628 766 13624 823
rect 5504 756 13624 766
rect 13457 727 13624 756
rect 2349 717 13377 727
rect 2349 713 13220 717
rect 5549 657 5835 713
rect 9035 657 9321 713
rect 12521 657 13220 713
rect 2349 647 13377 657
rect 13457 717 16735 727
rect 13614 714 16578 717
rect 13614 657 14296 714
rect 15896 657 16578 714
rect 13457 647 16735 657
rect 5553 609 5609 619
rect 5553 399 5609 409
rect 12525 609 12581 619
rect 12525 399 12581 409
rect 2349 361 13377 371
rect 5549 305 5835 361
rect 9035 305 9321 361
rect 12521 305 13220 361
rect 2349 301 13220 305
rect 2349 291 13377 301
rect 13457 361 16735 371
rect 13614 304 14296 361
rect 15896 304 16578 361
rect 13614 301 16578 304
rect 13457 291 16735 301
rect 2349 185 13377 195
rect 2349 181 13220 185
rect 5549 125 5835 181
rect 9035 125 9321 181
rect 12521 125 13220 181
rect 2349 115 13377 125
rect 13457 185 16735 195
rect 13614 182 16578 185
rect 13614 125 14296 182
rect 15896 125 16578 182
rect 13457 115 16735 125
rect 5553 77 5609 87
rect 5553 -133 5609 -123
rect 12525 77 12581 87
rect 12525 -133 12581 -123
rect 15902 77 16974 87
rect 15954 76 16974 77
rect 15954 -123 16822 76
rect 15902 -124 16822 -123
rect 16963 -124 16974 76
rect 15902 -133 16974 -124
rect 2349 -171 13377 -161
rect 5549 -227 5835 -171
rect 9035 -227 9321 -171
rect 12521 -227 13220 -171
rect 2349 -231 13220 -227
rect 2349 -241 13377 -231
rect 13457 -171 16735 -161
rect 13614 -228 14296 -171
rect 15896 -228 16577 -171
rect 13614 -231 16577 -228
rect 16734 -231 16735 -171
rect 13457 -241 16735 -231
rect 5504 -279 13614 -269
rect 5661 -339 12471 -279
rect 12628 -339 13457 -279
rect 5504 -349 13614 -339
<< via2 >>
rect 13457 1721 13614 1781
rect 16578 1721 16735 1781
rect 16823 1473 16964 1673
rect 13457 1365 13614 1425
rect 16578 1365 16735 1425
rect 13457 1189 13614 1249
rect 16578 1189 16735 1249
rect 13457 833 13614 893
rect 16578 833 16735 893
rect 5504 766 5661 826
rect 12471 766 12628 826
rect 13220 657 13377 717
rect 13457 657 13614 717
rect 16578 657 16735 717
rect 5553 409 5555 609
rect 5555 409 5607 609
rect 5607 409 5609 609
rect 12525 409 12527 609
rect 12527 409 12579 609
rect 12579 409 12581 609
rect 13220 301 13377 361
rect 13457 301 13614 361
rect 16578 301 16735 361
rect 13220 125 13377 185
rect 13457 125 13614 185
rect 16578 125 16735 185
rect 5553 -123 5555 77
rect 5555 -123 5607 77
rect 5607 -123 5609 77
rect 12525 -123 12527 77
rect 12527 -123 12579 77
rect 12579 -123 12581 77
rect 16822 -124 16963 76
rect 13220 -231 13377 -171
rect 13457 -231 13614 -171
rect 16577 -231 16734 -171
rect 5504 -339 5661 -279
rect 12471 -339 12628 -279
rect 13457 -339 13614 -279
<< metal3 >>
rect 13447 1781 13624 1792
rect 13447 1721 13457 1781
rect 13614 1721 13624 1781
rect 13447 1425 13624 1721
rect 13447 1365 13457 1425
rect 13614 1365 13624 1425
rect 13447 1249 13624 1365
rect 13447 1189 13457 1249
rect 13614 1189 13624 1249
rect 13447 893 13624 1189
rect 13447 833 13457 893
rect 13614 833 13624 893
rect 5494 826 5671 831
rect 5494 766 5504 826
rect 5661 766 5671 826
rect 5494 761 5671 766
rect 12461 826 12638 831
rect 12461 766 12471 826
rect 12628 766 12638 826
rect 12461 761 12638 766
rect 5543 609 5619 761
rect 5543 409 5553 609
rect 5609 409 5619 609
rect 5543 77 5619 409
rect 5543 -123 5553 77
rect 5609 -123 5619 77
rect 5543 -274 5619 -123
rect 12515 609 12591 761
rect 12515 409 12525 609
rect 12581 409 12591 609
rect 12515 77 12591 409
rect 12515 -123 12525 77
rect 12581 -123 12591 77
rect 12515 -274 12591 -123
rect 13210 717 13387 728
rect 13210 657 13220 717
rect 13377 657 13387 717
rect 13210 361 13387 657
rect 13210 301 13220 361
rect 13377 301 13387 361
rect 13210 185 13387 301
rect 13210 125 13220 185
rect 13377 125 13387 185
rect 13210 -171 13387 125
rect 13210 -231 13220 -171
rect 13377 -231 13387 -171
rect 13210 -236 13387 -231
rect 13447 717 13624 833
rect 13447 657 13457 717
rect 13614 657 13624 717
rect 13447 361 13624 657
rect 13447 301 13457 361
rect 13614 301 13624 361
rect 13447 185 13624 301
rect 13447 125 13457 185
rect 13614 125 13624 185
rect 13447 -171 13624 125
rect 13447 -231 13457 -171
rect 13614 -231 13624 -171
rect 5494 -279 5671 -274
rect 5494 -339 5504 -279
rect 5661 -339 5671 -279
rect 5494 -344 5671 -339
rect 12461 -279 12638 -274
rect 12461 -339 12471 -279
rect 12628 -339 12638 -279
rect 12461 -344 12638 -339
rect 13447 -279 13624 -231
rect 16567 1781 16745 1791
rect 16567 1721 16578 1781
rect 16735 1721 16745 1781
rect 16567 1425 16745 1721
rect 16567 1365 16578 1425
rect 16735 1365 16745 1425
rect 16567 1249 16745 1365
rect 16567 1189 16578 1249
rect 16735 1189 16745 1249
rect 16567 893 16745 1189
rect 16567 833 16578 893
rect 16735 833 16745 893
rect 16567 717 16745 833
rect 16567 657 16578 717
rect 16735 657 16745 717
rect 16567 361 16745 657
rect 16567 301 16578 361
rect 16735 301 16745 361
rect 16567 185 16745 301
rect 16567 125 16578 185
rect 16735 125 16745 185
rect 16567 -171 16745 125
rect 16567 -231 16577 -171
rect 16734 -231 16745 -171
rect 16567 -241 16745 -231
rect 16805 1673 16974 1683
rect 16805 1473 16823 1673
rect 16964 1473 16974 1673
rect 16805 76 16974 1473
rect 16805 -124 16822 76
rect 16963 -124 16974 76
rect 16805 -236 16974 -124
rect 13447 -339 13457 -279
rect 13614 -339 13624 -279
rect 13447 -375 13624 -339
use trans_gate  x1
timestamp 1712344797
transform 1 0 -674 0 1 -2250
box 0 -2052 3413 715
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[0]
timestamp 1712597941
transform 1 0 11537 0 1 -2072
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[1]
timestamp 1712597941
transform 1 0 11537 0 1 -3364
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[0]
timestamp 1712597941
transform 1 0 11537 0 1 -2718
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[1]
timestamp 1712597941
transform 1 0 11537 0 1 -4010
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[0]
timestamp 1712343889
transform 1 0 15096 0 1 1041
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[1]
timestamp 1712343889
transform 1 0 15096 0 1 509
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM4[0]
timestamp 1712669456
transform 1 0 7435 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1712671997
transform 1 0 7435 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[0]
timestamp 1712343889
transform 1 0 15096 0 1 1573
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[1]
timestamp 1712343889
transform 1 0 15096 0 1 -23
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[0]
timestamp 1712669456
transform 1 0 3949 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1712671997
transform 1 0 3949 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[2]
timestamp 1712669456
transform 1 0 10921 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1712671997
transform 1 0 10921 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1712343889
transform 1 0 14601 0 1 -1841
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_697RXD  XM8
timestamp 1712343889
transform 1 0 14601 0 1 -2906
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1712343889
transform 1 0 16150 0 1 -1649
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1712343889
transform 1 0 16050 0 1 -3126
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1712343889
transform 1 0 7247 0 1 -2114
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1712343889
transform 1 0 7485 0 1 -1380
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1712343889
transform 1 0 8947 0 1 -2895
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1712343889
transform 1 0 8939 0 1 -3612
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1712343889
transform 1 0 12397 0 1 2117
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1712343889
transform 1 0 11109 0 1 2136
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1712343889
transform 1 0 14131 0 1 -3659
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1712343889
transform 1 0 4155 0 1 -1447
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1712343889
transform 1 0 4155 0 1 -2201
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[0]
timestamp 1712671997
transform 1 0 13910 0 1 2105
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[1]
timestamp 1712671997
transform 1 0 13910 0 1 1573
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[2]
timestamp 1712671997
transform 1 0 13910 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[3]
timestamp 1712671997
transform 1 0 13910 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712671997
transform 1 0 13910 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712671997
transform 1 0 13910 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712671997
transform 1 0 16282 0 1 2105
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712671997
transform 1 0 16282 0 1 1573
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712671997
transform 1 0 16282 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712671997
transform 1 0 16282 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712671997
transform 1 0 16282 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712671997
transform 1 0 16282 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712671997
transform 1 0 1963 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712671997
transform 1 0 1963 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712671997
transform 1 0 1963 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712671997
transform 1 0 1963 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[16]
timestamp 1712671997
transform 1 0 12907 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[17]
timestamp 1712671997
transform 1 0 12907 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[18]
timestamp 1712671997
transform 1 0 12907 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[19]
timestamp 1712671997
transform 1 0 12907 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[0]
timestamp 1712343889
transform 1 0 15096 0 1 2105
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[1]
timestamp 1712343889
transform 1 0 15096 0 1 -555
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712671997
transform 1 0 3949 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712671997
transform 1 0 7435 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712671997
transform 1 0 10921 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712671997
transform 1 0 3949 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712671997
transform 1 0 7435 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712671997
transform 1 0 10921 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712600458
transform 1 0 10199 0 1 -1456
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712600458
transform 1 0 10199 0 1 -4626
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712600458
transform 1 0 12875 0 1 -1456
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712600458
transform 1 0 12875 0 1 -4626
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712599722
transform 1 0 11537 0 1 -1456
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712599722
transform 1 0 11537 0 1 -4626
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712597941
transform 1 0 10199 0 1 -2072
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712597941
transform 1 0 10199 0 1 -2718
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712597941
transform 1 0 10199 0 1 -3364
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712597941
transform 1 0 10199 0 1 -4010
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[4]
timestamp 1712597941
transform 1 0 12875 0 1 -2072
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[5]
timestamp 1712597941
transform 1 0 12875 0 1 -2718
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[6]
timestamp 1712597941
transform 1 0 12875 0 1 -3364
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[7]
timestamp 1712597941
transform 1 0 12875 0 1 -4010
box -328 -388 328 388
<< labels >>
flabel metal1 20126 -2729 20326 -2529 0 FreeSans 256 180 0 0 dvdd
port 0 nsew
flabel metal1 20126 -2329 20326 -2129 0 FreeSans 256 180 0 0 out
port 1 nsew
flabel metal1 20126 -329 20326 -129 0 FreeSans 256 180 0 0 vss
port 6 nsew
flabel metal1 20126 -729 20326 -529 0 FreeSans 256 180 0 0 ibias
port 5 nsew
flabel metal1 20126 -1129 20326 -929 0 FreeSans 256 180 0 0 ena
port 4 nsew
flabel metal1 20126 -1529 20326 -1329 0 FreeSans 256 180 0 0 vin
port 3 nsew
flabel metal1 20126 -1929 20326 -1729 0 FreeSans 256 180 0 0 vref
port 2 nsew
<< end >>

* NGSPICE file created from sky130_vbl_ip__overvoltage.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_LV9PDH a_8742_125# a_n3732_n557# a_1560_125#
+ a_3828_n557# a_n7512_n557# a_804_n557# a_7608_n557# a_n4110_n557# a_3072_125# a_4206_n557#
+ a_4584_125# a_n4110_125# a_6096_125# a_n5622_125# a_6852_n557# a_n4866_n557# a_n1464_n557#
+ a_3450_n557# a_48_125# a_n8646_n557# a_7230_n557# a_n5244_n557# a_n7134_125# a_n8646_125#
+ a_n1464_125# a_n9024_n557# a_n2976_125# a_804_125# a_2316_125# a_3828_125# a_n7890_n557#
+ a_5340_125# a_7986_n557# a_n4488_125# a_4584_n557# a_n2598_n557# a_1182_n557# a_6852_125#
+ a_8364_n557# a_n6378_n557# a_8364_125# a_1182_125# a_2694_125# a_n2220_125# a_n1842_n557#
+ a_48_n557# a_1938_n557# a_n3732_125# a_n708_125# a_n5622_n557# a_n2220_n557# a_5718_n557#
+ a_2316_n557# a_6096_n557# a_n5244_125# a_n6000_n557# a_n6756_125# a_7608_125# a_n8268_125#
+ a_n2976_n557# a_4962_n557# a_n1086_125# a_1560_n557# a_1938_125# a_n2598_125# a_3450_125#
+ a_4962_125# a_8742_n557# a_5340_n557# a_n6756_n557# a_426_125# a_n3354_n557# a_6474_125#
+ a_n7134_n557# a_426_n557# a_7986_125# a_n708_n557# a_n6000_125# a_n7512_125# a_2694_n557#
+ a_n1842_125# a_6474_n557# a_3072_n557# a_n4488_n557# a_n1086_n557# a_n330_125# a_n9024_125#
+ a_n3354_125# a_n8268_n557# a_n4866_125# a_n330_n557# a_n7890_125# a_4206_125# a_5718_125#
+ a_7230_125# 0 a_n6378_125#
X0 a_n8646_125# a_n8646_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X1 a_n6000_125# a_n6000_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X2 a_n1464_125# a_n1464_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X3 a_6474_125# a_6474_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X4 a_804_125# a_804_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X5 a_n7134_125# a_n7134_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X6 a_n4488_125# a_n4488_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X7 a_5718_125# a_5718_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X8 a_n1842_125# a_n1842_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X9 a_6852_125# a_6852_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X10 a_n7512_125# a_n7512_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X11 a_n4866_125# a_n4866_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X12 a_4206_125# a_4206_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X13 a_5340_125# a_5340_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X14 a_n330_125# a_n330_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X15 a_2694_125# a_2694_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X16 a_n7890_125# a_n7890_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X17 a_n3354_125# a_n3354_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X18 a_n2220_125# a_n2220_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X19 a_8364_125# a_8364_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X20 a_1182_125# a_1182_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X21 a_1938_125# a_1938_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X22 a_n9024_125# a_n9024_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X23 a_n708_125# a_n708_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X24 a_48_125# a_48_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X25 a_n6378_125# a_n6378_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X26 a_n3732_125# a_n3732_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X27 a_7608_125# a_7608_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X28 a_8742_125# a_8742_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X29 a_1560_125# a_1560_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X30 a_n6756_125# a_n6756_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X31 a_7230_125# a_7230_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X32 a_4584_125# a_4584_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X33 a_n5244_125# a_n5244_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X34 a_n4110_125# a_n4110_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X35 a_n2598_125# a_n2598_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X36 a_3072_125# a_3072_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X37 a_3828_125# a_3828_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X38 a_4962_125# a_4962_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X39 a_n8268_125# a_n8268_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X40 a_n5622_125# a_n5622_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X41 a_n2976_125# a_n2976_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X42 a_n1086_125# a_n1086_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X43 a_6096_125# a_6096_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X44 a_7986_125# a_7986_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X45 a_426_125# a_426_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X46 a_2316_125# a_2316_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X47 a_3450_125# a_3450_n557# 0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
C0 a_n7512_125# a_n7512_n557# 0.063641f
C1 a_5718_125# a_6096_125# 0.296258f
C2 a_n1464_125# a_n1086_125# 0.296258f
C3 a_n8646_125# a_n9024_125# 0.296258f
C4 a_3072_125# a_2694_125# 0.296258f
C5 a_1560_n557# a_1938_n557# 0.296258f
C6 a_7986_n557# a_7986_125# 0.063641f
C7 a_n4110_125# a_n3732_125# 0.296258f
C8 a_n5244_125# a_n5622_125# 0.296258f
C9 a_7986_n557# a_7608_n557# 0.296258f
C10 a_8742_n557# a_8742_125# 0.063641f
C11 a_3828_125# a_3828_n557# 0.063641f
C12 a_804_n557# a_426_n557# 0.296258f
C13 a_6852_n557# a_6474_n557# 0.296258f
C14 a_8364_125# a_8742_125# 0.296258f
C15 a_4206_n557# a_3828_n557# 0.296258f
C16 a_n8268_n557# a_n7890_n557# 0.296258f
C17 a_1560_125# a_1938_125# 0.296258f
C18 a_n2598_n557# a_n2976_n557# 0.296258f
C19 a_7230_125# a_6852_125# 0.296258f
C20 a_1182_125# a_1182_n557# 0.063641f
C21 a_7230_n557# a_6852_n557# 0.296258f
C22 a_n6756_n557# a_n6756_125# 0.063641f
C23 a_n2220_125# a_n2598_125# 0.296258f
C24 a_n6378_125# a_n6378_n557# 0.063641f
C25 a_804_n557# a_804_125# 0.063641f
C26 a_7986_n557# a_8364_n557# 0.296258f
C27 a_4584_125# a_4584_n557# 0.063641f
C28 a_n4866_125# a_n4488_125# 0.296258f
C29 a_1182_n557# a_1560_n557# 0.296258f
C30 a_n330_n557# a_48_n557# 0.296258f
C31 a_7608_125# a_7230_125# 0.296258f
C32 a_n708_n557# a_n330_n557# 0.296258f
C33 a_2316_125# a_2694_125# 0.296258f
C34 a_3072_125# a_3072_n557# 0.063641f
C35 a_6474_125# a_6474_n557# 0.063641f
C36 a_n8646_n557# a_n9024_n557# 0.296258f
C37 a_7608_125# a_7986_125# 0.296258f
C38 a_n3354_n557# a_n3732_n557# 0.296258f
C39 a_n330_125# a_48_125# 0.296258f
C40 a_n1086_125# a_n708_125# 0.296258f
C41 a_2316_n557# a_2316_125# 0.063641f
C42 a_4206_125# a_3828_125# 0.296258f
C43 a_n2220_125# a_n1842_125# 0.296258f
C44 a_n7134_125# a_n6756_125# 0.296258f
C45 a_3072_125# a_3450_125# 0.296258f
C46 a_n2976_125# a_n2976_n557# 0.063641f
C47 a_n5244_n557# a_n4866_n557# 0.296258f
C48 a_n2976_125# a_n3354_125# 0.296258f
C49 a_n708_n557# a_n1086_n557# 0.296258f
C50 a_7608_n557# a_7608_125# 0.063641f
C51 a_4206_n557# a_4206_125# 0.063641f
C52 a_n3732_n557# a_n3732_125# 0.063641f
C53 a_3828_125# a_3450_125# 0.296258f
C54 a_6096_125# a_6096_n557# 0.063641f
C55 a_n8268_125# a_n8268_n557# 0.063641f
C56 a_n8268_n557# a_n8646_n557# 0.296258f
C57 a_n2598_n557# a_n2220_n557# 0.296258f
C58 a_5718_125# a_5340_125# 0.296258f
C59 a_n1464_n557# a_n1842_n557# 0.296258f
C60 a_n330_125# a_n708_125# 0.296258f
C61 a_1938_125# a_1938_n557# 0.063641f
C62 a_n5622_125# a_n6000_125# 0.296258f
C63 a_n4110_125# a_n4110_n557# 0.063641f
C64 a_n5622_n557# a_n5622_125# 0.063641f
C65 a_n8268_125# a_n8646_125# 0.296258f
C66 a_48_n557# a_426_n557# 0.296258f
C67 a_n8646_n557# a_n8646_125# 0.063641f
C68 a_n4110_n557# a_n4488_n557# 0.296258f
C69 a_n6000_n557# a_n6000_125# 0.063641f
C70 a_5340_125# a_5340_n557# 0.063641f
C71 a_4962_125# a_5340_125# 0.296258f
C72 a_n5622_n557# a_n6000_n557# 0.296258f
C73 a_5718_125# a_5718_n557# 0.063641f
C74 a_426_125# a_426_n557# 0.063641f
C75 a_n1464_125# a_n1842_125# 0.296258f
C76 a_2694_n557# a_2694_125# 0.063641f
C77 a_4962_125# a_4584_125# 0.296258f
C78 a_5718_n557# a_5340_n557# 0.296258f
C79 a_n5244_n557# a_n5244_125# 0.063641f
C80 a_n1842_n557# a_n2220_n557# 0.296258f
C81 a_n6756_n557# a_n7134_n557# 0.296258f
C82 a_426_125# a_804_125# 0.296258f
C83 a_2694_n557# a_2316_n557# 0.296258f
C84 a_n4110_125# a_n4488_125# 0.296258f
C85 a_1182_n557# a_804_n557# 0.296258f
C86 a_n4866_125# a_n4866_n557# 0.063641f
C87 a_8364_125# a_7986_125# 0.296258f
C88 a_3450_n557# a_3828_n557# 0.296258f
C89 a_n4488_125# a_n4488_n557# 0.063641f
C90 a_4962_n557# a_4584_n557# 0.296258f
C91 a_6852_n557# a_6852_125# 0.063641f
C92 a_n2598_n557# a_n2598_125# 0.063641f
C93 a_4206_n557# a_4584_n557# 0.296258f
C94 a_n7134_125# a_n7134_n557# 0.063641f
C95 a_n7890_125# a_n7890_n557# 0.063641f
C96 a_n6756_n557# a_n6378_n557# 0.296258f
C97 a_n1464_n557# a_n1086_n557# 0.296258f
C98 a_7230_n557# a_7230_125# 0.063641f
C99 a_n3732_n557# a_n4110_n557# 0.296258f
C100 a_n6756_125# a_n6378_125# 0.296258f
C101 a_1182_125# a_1560_125# 0.296258f
C102 a_8742_n557# a_8364_n557# 0.296258f
C103 a_2694_n557# a_3072_n557# 0.296258f
C104 a_8364_125# a_8364_n557# 0.063641f
C105 a_1560_125# a_1560_n557# 0.063641f
C106 a_48_125# a_48_n557# 0.063641f
C107 a_6096_125# a_6474_125# 0.296258f
C108 a_n330_125# a_n330_n557# 0.063641f
C109 a_n1086_125# a_n1086_n557# 0.063641f
C110 a_n5244_125# a_n4866_125# 0.296258f
C111 a_3450_n557# a_3072_n557# 0.296258f
C112 a_n7512_n557# a_n7134_n557# 0.296258f
C113 a_2316_n557# a_1938_n557# 0.296258f
C114 a_48_125# a_426_125# 0.296258f
C115 a_n3354_n557# a_n2976_n557# 0.296258f
C116 a_n3354_n557# a_n3354_125# 0.063641f
C117 a_n6000_n557# a_n6378_n557# 0.296258f
C118 a_7608_n557# a_7230_n557# 0.296258f
C119 a_6474_125# a_6852_125# 0.296258f
C120 a_n7512_n557# a_n7890_n557# 0.296258f
C121 a_1182_125# a_804_125# 0.296258f
C122 a_3450_n557# a_3450_125# 0.063641f
C123 a_n7890_125# a_n7512_125# 0.296258f
C124 a_5718_n557# a_6096_n557# 0.296258f
C125 a_n2976_125# a_n2598_125# 0.296258f
C126 a_n3354_125# a_n3732_125# 0.296258f
C127 a_n9024_n557# a_n9024_125# 0.063641f
C128 a_n6378_125# a_n6000_125# 0.296258f
C129 a_n7512_125# a_n7134_125# 0.296258f
C130 a_n708_n557# a_n708_125# 0.063641f
C131 a_4584_125# a_4206_125# 0.296258f
C132 a_n5244_n557# a_n5622_n557# 0.296258f
C133 a_6096_n557# a_6474_n557# 0.296258f
C134 a_4962_n557# a_5340_n557# 0.296258f
C135 a_4962_125# a_4962_n557# 0.063641f
C136 a_n2220_125# a_n2220_n557# 0.063641f
C137 a_n8268_125# a_n7890_125# 0.296258f
C138 a_n1464_n557# a_n1464_125# 0.063641f
C139 a_n4866_n557# a_n4488_n557# 0.296258f
C140 a_n1842_n557# a_n1842_125# 0.063641f
C141 a_1938_125# a_2316_125# 0.296258f
C142 a_8742_n557# 0 0.562823f
C143 a_8742_125# 0 0.562823f
C144 a_8364_n557# 0 0.354294f
C145 a_8364_125# 0 0.354294f
C146 a_7986_n557# 0 0.354294f
C147 a_7986_125# 0 0.354294f
C148 a_7608_n557# 0 0.354294f
C149 a_7608_125# 0 0.354294f
C150 a_7230_n557# 0 0.354294f
C151 a_7230_125# 0 0.354294f
C152 a_6852_n557# 0 0.354294f
C153 a_6852_125# 0 0.354294f
C154 a_6474_n557# 0 0.354294f
C155 a_6474_125# 0 0.354294f
C156 a_6096_n557# 0 0.354294f
C157 a_6096_125# 0 0.354294f
C158 a_5718_n557# 0 0.354294f
C159 a_5718_125# 0 0.354294f
C160 a_5340_n557# 0 0.354294f
C161 a_5340_125# 0 0.354294f
C162 a_4962_n557# 0 0.354294f
C163 a_4962_125# 0 0.354294f
C164 a_4584_n557# 0 0.354294f
C165 a_4584_125# 0 0.354294f
C166 a_4206_n557# 0 0.354294f
C167 a_4206_125# 0 0.354294f
C168 a_3828_n557# 0 0.354294f
C169 a_3828_125# 0 0.354294f
C170 a_3450_n557# 0 0.354294f
C171 a_3450_125# 0 0.354294f
C172 a_3072_n557# 0 0.354294f
C173 a_3072_125# 0 0.354294f
C174 a_2694_n557# 0 0.354294f
C175 a_2694_125# 0 0.354294f
C176 a_2316_n557# 0 0.354294f
C177 a_2316_125# 0 0.354294f
C178 a_1938_n557# 0 0.354294f
C179 a_1938_125# 0 0.354294f
C180 a_1560_n557# 0 0.354294f
C181 a_1560_125# 0 0.354294f
C182 a_1182_n557# 0 0.354294f
C183 a_1182_125# 0 0.354294f
C184 a_804_n557# 0 0.354294f
C185 a_804_125# 0 0.354294f
C186 a_426_n557# 0 0.354294f
C187 a_426_125# 0 0.354294f
C188 a_48_n557# 0 0.354294f
C189 a_48_125# 0 0.354294f
C190 a_n330_n557# 0 0.354294f
C191 a_n330_125# 0 0.354294f
C192 a_n708_n557# 0 0.354294f
C193 a_n708_125# 0 0.354294f
C194 a_n1086_n557# 0 0.354294f
C195 a_n1086_125# 0 0.354294f
C196 a_n1464_n557# 0 0.354294f
C197 a_n1464_125# 0 0.354294f
C198 a_n1842_n557# 0 0.354294f
C199 a_n1842_125# 0 0.354294f
C200 a_n2220_n557# 0 0.354294f
C201 a_n2220_125# 0 0.354294f
C202 a_n2598_n557# 0 0.354294f
C203 a_n2598_125# 0 0.354294f
C204 a_n2976_n557# 0 0.354294f
C205 a_n2976_125# 0 0.354294f
C206 a_n3354_n557# 0 0.354294f
C207 a_n3354_125# 0 0.354294f
C208 a_n3732_n557# 0 0.354294f
C209 a_n3732_125# 0 0.354294f
C210 a_n4110_n557# 0 0.354294f
C211 a_n4110_125# 0 0.354294f
C212 a_n4488_n557# 0 0.354294f
C213 a_n4488_125# 0 0.354294f
C214 a_n4866_n557# 0 0.354294f
C215 a_n4866_125# 0 0.354294f
C216 a_n5244_n557# 0 0.354294f
C217 a_n5244_125# 0 0.354294f
C218 a_n5622_n557# 0 0.354294f
C219 a_n5622_125# 0 0.354294f
C220 a_n6000_n557# 0 0.354294f
C221 a_n6000_125# 0 0.354294f
C222 a_n6378_n557# 0 0.354294f
C223 a_n6378_125# 0 0.354294f
C224 a_n6756_n557# 0 0.354294f
C225 a_n6756_125# 0 0.354294f
C226 a_n7134_n557# 0 0.354294f
C227 a_n7134_125# 0 0.354294f
C228 a_n7512_n557# 0 0.354294f
C229 a_n7512_125# 0 0.354294f
C230 a_n7890_n557# 0 0.354294f
C231 a_n7890_125# 0 0.354294f
C232 a_n8268_n557# 0 0.354294f
C233 a_n8268_125# 0 0.354294f
C234 a_n8646_n557# 0 0.354294f
C235 a_n8646_125# 0 0.354294f
C236 a_n9024_n557# 0 0.562823f
C237 a_n9024_125# 0 0.562823f
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_H3F4MM a_1182_1930# a_n4488_n1826# a_7986_n1826#
+ a_n6378_n2362# a_n7890_5150# a_n7890_n5582# a_7986_5150# a_4584_5150# a_n2598_5150#
+ a_1182_5150# a_8364_1930# a_n6378_1930# a_n4866_n1826# a_n6756_n2362# a_8364_5150#
+ a_n6378_5150# a_n2598_n1826# a_n6000_n5582# a_n4488_n2362# a_n3732_1394# a_7986_n2362#
+ a_3828_1394# a_426_n5582# a_7230_n5582# a_7608_n5582# a_n2976_n1826# a_n4866_n2362#
+ a_n7512_1394# a_n4110_1394# a_804_1394# a_7608_1394# a_4206_1394# a_4206_n1826#
+ a_n1842_1930# a_n4110_n5582# a_804_n5582# a_n2598_n2362# a_48_1930# a_1938_1930#
+ a_5340_n5582# a_n1842_5150# a_5718_n5582# a_48_5150# a_1938_5150# a_n5622_1930#
+ a_n2976_n2362# a_n2220_1930# a_5718_1930# a_3072_n5582# a_2316_1930# a_n9024_n1826#
+ a_6096_1930# a_2316_n1826# a_4206_n2362# a_n2220_n5582# a_n5622_5150# a_n2220_5150#
+ a_5718_5150# a_2316_5150# a_6852_1394# a_n6000_1930# a_6096_5150# a_n4866_1394#
+ a_3450_1394# a_3450_n5582# a_3828_n5582# a_n1464_1394# a_n8268_n5582# a_n6000_5150#
+ a_1182_n5582# a_n7134_n1826# a_n9024_n2362# a_2316_n2362# a_n8646_1394# a_7230_1394#
+ a_n5244_1394# a_8364_n1826# a_4962_1930# a_n2976_1930# a_1560_1930# a_n8646_n5582#
+ a_1560_n5582# a_n7512_n1826# a_1938_n5582# a_6096_n1826# a_n9024_1394# a_4962_5150#
+ a_n2976_5150# a_n6378_n5582# a_n5244_n1826# a_n7134_n2362# a_1560_5150# a_8742_n1826#
+ a_8742_1930# a_n6756_1930# a_5340_1930# a_n3354_1930# a_n330_n1826# a_6474_n1826#
+ a_n708_n1826# a_8364_n2362# a_8742_5150# a_n6756_n5582# a_n6756_5150# a_n5622_n1826#
+ a_5340_5150# a_n7512_n2362# a_48_n1826# a_n7890_1394# a_n3354_5150# a_6096_n2362#
+ a_n7134_1930# a_7986_1394# a_n4488_n5582# a_426_1930# a_4584_1394# a_7986_n5582#
+ a_n3354_n1826# a_n2598_1394# a_6852_n1826# a_n5244_n2362# a_8742_n2362# a_1182_1394#
+ a_n708_1930# a_n7134_5150# a_n1086_n1826# a_426_5150# a_4584_n1826# a_n330_n2362#
+ a_6474_n2362# a_n708_n2362# a_8364_1394# a_n4866_n5582# a_n3732_n1826# a_n6378_1394#
+ a_n5622_n2362# a_48_n2362# a_n708_5150# a_2694_1930# a_n2598_n5582# a_n1464_n1826#
+ a_4962_n1826# a_n3354_n2362# a_6852_n2362# a_2694_5150# a_2694_n1826# a_n1086_n2362#
+ a_4584_n2362# a_6474_1930# a_n2976_n5582# a_n4488_1930# a_n1842_n1826# a_n3732_n2362#
+ a_3072_1930# a_n1086_1930# a_4206_n5582# a_6474_5150# a_n1464_n2362# a_4962_n2362#
+ a_n4488_5150# a_3072_5150# a_n1842_1394# a_n1086_5150# a_n8268_1930# a_48_1394#
+ a_1938_1394# a_2694_n2362# a_n330_1930# a_n1842_n2362# a_n8268_5150# a_n5622_1394#
+ a_n9024_n5582# a_n2220_1394# a_2316_n5582# a_5718_1394# a_n7890_n1826# a_n330_5150#
+ a_2316_1394# a_6096_1394# a_n6000_1394# a_n3732_1930# a_n7134_n5582# a_3828_1930#
+ a_n6000_n1826# a_n7890_n2362# a_n3732_5150# a_8364_n5582# a_426_n1826# a_7230_n1826#
+ a_3828_5150# a_7608_n1826# a_n7512_1930# a_n7512_n5582# a_n4110_1930# a_804_1930#
+ a_7608_1930# a_4962_1394# a_n2976_1394# a_4206_1930# a_1560_1394# a_6096_n5582#
+ a_n7512_5150# a_n5244_n5582# a_n4110_n1826# a_8742_n5582# a_804_n1826# a_n6000_n2362#
+ a_n4110_5150# a_804_5150# a_7608_5150# a_4206_5150# a_8742_1394# a_n6756_1394# a_5340_1394#
+ a_n3354_1394# a_6474_n5582# a_n330_n5582# a_n708_n5582# a_5340_n1826# a_426_n2362#
+ a_5718_n1826# a_7230_n2362# a_7608_n2362# a_n5622_n5582# a_48_n5582# a_3072_n1826#
+ a_n7134_1394# a_n3354_n5582# a_6852_n5582# a_n2220_n1826# a_n4110_n2362# a_804_n2362#
+ a_426_1394# a_6852_1930# a_n4866_1930# a_3450_1930# a_n1464_1930# a_n1086_n5582#
+ a_4584_n5582# a_n708_1394# a_3450_n1826# a_5340_n2362# a_3828_n1826# a_5718_n2362#
+ a_n3732_n5582# a_6852_5150# a_n4866_5150# a_3450_5150# a_n1464_5150# a_n8268_n1826#
+ a_1182_n1826# a_n8646_1930# a_3072_n2362# a_7230_1930# a_n5244_1930# a_n1464_n5582#
+ a_4962_n5582# a_n2220_n2362# a_2694_1394# a_n8646_5150# a_7230_5150# a_2694_n5582#
+ a_n8646_n1826# a_n5244_5150# a_1560_n1826# a_1938_n1826# a_3450_n2362# a_3828_n2362#
+ a_n9024_1930# a_n1842_n5582# a_6474_1394# a_n4488_1394# a_3072_1394# a_n6378_n1826#
+ a_n8268_n2362# a_n1086_1394# a_1182_n2362# a_n9024_5150# a_n8268_1394# a_n7890_1930#
+ a_n6756_n1826# a_n8646_n2362# a_1560_n2362# a_1938_n2362# a_7986_1930# 0 a_4584_1930#
+ a_n2598_1930# a_n330_1394#
X0 a_n1464_n2362# a_n1464_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X1 a_n3732_n2362# a_n3732_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X2 a_426_n2362# a_426_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X3 a_n4110_5150# a_n4110_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X4 a_n5244_5150# a_n5244_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X5 a_n2598_5150# a_n2598_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X6 a_3072_5150# a_3072_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X7 a_3828_5150# a_3828_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X8 a_4962_5150# a_4962_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X9 a_n9024_1394# a_n9024_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X10 a_6474_1394# a_6474_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X11 a_n8268_5150# a_n8268_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X12 a_8742_1394# a_8742_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X13 a_5718_1394# a_5718_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X14 a_n330_1394# a_n330_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X15 a_n9024_n2362# a_n9024_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X16 a_3072_1394# a_3072_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X17 a_n7890_1394# a_n7890_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X18 a_n5622_5150# a_n5622_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X19 a_5340_1394# a_5340_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X20 a_2316_1394# a_2316_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X21 a_n1086_5150# a_n1086_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X22 a_6096_5150# a_6096_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X23 a_6474_n2362# a_6474_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X24 a_8742_n2362# a_8742_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X25 a_5718_n2362# a_5718_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X26 a_n330_n2362# a_n330_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X27 a_7986_5150# a_7986_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X28 a_n4488_1394# a_n4488_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X29 a_n2976_5150# a_n2976_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X30 a_2316_5150# a_2316_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X31 a_n6756_1394# a_n6756_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X32 a_426_5150# a_426_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X33 a_3450_5150# a_3450_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X34 a_3072_n2362# a_3072_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X35 a_n7890_n2362# a_n7890_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X36 a_5340_n2362# a_5340_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X37 a_2316_n2362# a_2316_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X38 a_n1086_1394# a_n1086_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X39 a_n3354_1394# a_n3354_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X40 a_n4488_n2362# a_n4488_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X41 a_n5622_1394# a_n5622_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X42 a_n6756_n2362# a_n6756_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X43 a_n1086_n2362# a_n1086_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X44 a_n8646_5150# a_n8646_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X45 a_n3354_n2362# a_n3354_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X46 a_n5622_n2362# a_n5622_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X47 a_n6000_5150# a_n6000_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X48 a_6474_5150# a_6474_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X49 a_n1464_5150# a_n1464_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X50 a_804_5150# a_804_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X51 a_n7134_5150# a_n7134_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X52 a_6096_1394# a_6096_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X53 a_n4488_5150# a_n4488_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X54 a_8364_1394# a_8364_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X55 a_7608_1394# a_7608_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X56 a_n1842_5150# a_n1842_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X57 a_5718_5150# a_5718_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X58 a_6852_5150# a_6852_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X59 a_6096_n2362# a_6096_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X60 a_7230_1394# a_7230_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X61 a_4206_1394# a_4206_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X62 a_8364_n2362# a_8364_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X63 a_7608_n2362# a_7608_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X64 a_n6378_1394# a_n6378_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X65 a_n8646_1394# a_n8646_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X66 a_7230_n2362# a_7230_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X67 a_4206_n2362# a_4206_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X68 a_n2220_1394# a_n2220_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X69 a_n5244_1394# a_n5244_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X70 a_n6378_n2362# a_n6378_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X71 a_n7512_1394# a_n7512_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X72 a_n7512_5150# a_n7512_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X73 a_n8646_n2362# a_n8646_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X74 a_2694_1394# a_2694_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X75 a_n4866_5150# a_n4866_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X76 a_4206_5150# a_4206_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X77 a_4962_1394# a_4962_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X78 a_1938_1394# a_1938_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X79 a_5340_5150# a_5340_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X80 a_n2220_n2362# a_n2220_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X81 a_n5244_n2362# a_n5244_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X82 a_n7512_n2362# a_n7512_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X83 a_n330_5150# a_n330_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X84 a_2694_5150# a_2694_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X85 a_1560_1394# a_1560_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X86 a_2694_n2362# a_2694_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X87 a_4962_n2362# a_4962_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X88 a_1938_n2362# a_1938_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X89 a_48_1394# a_48_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X90 a_n2976_1394# a_n2976_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X91 a_1560_n2362# a_1560_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X92 a_48_n2362# a_48_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X93 a_n7890_5150# a_n7890_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X94 a_n1842_1394# a_n1842_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X95 a_n2220_5150# a_n2220_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X96 a_n2976_n2362# a_n2976_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X97 a_n3354_5150# a_n3354_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X98 a_8364_5150# a_8364_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X99 a_804_1394# a_804_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X100 a_1182_5150# a_1182_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X101 a_n1842_n2362# a_n1842_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X102 a_1938_5150# a_1938_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X103 a_804_n2362# a_804_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X104 a_n708_5150# a_n708_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X105 a_48_5150# a_48_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X106 a_n9024_5150# a_n9024_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X107 a_n8268_1394# a_n8268_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X108 a_n6378_5150# a_n6378_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X109 a_n3732_5150# a_n3732_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X110 a_7608_5150# a_7608_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X111 a_8742_5150# a_8742_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X112 a_7986_1394# a_7986_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X113 a_n4110_1394# a_n4110_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X114 a_n7134_1394# a_n7134_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X115 a_n8268_n2362# a_n8268_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X116 a_4584_1394# a_4584_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X117 a_1560_5150# a_1560_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X118 a_6852_1394# a_6852_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X119 a_3828_1394# a_3828_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X120 a_7986_n2362# a_7986_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X121 a_n4110_n2362# a_n4110_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X122 a_n7134_n2362# a_n7134_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X123 a_n708_1394# a_n708_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X124 a_1182_1394# a_1182_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X125 a_n6000_1394# a_n6000_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X126 a_3450_1394# a_3450_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X127 a_4584_n2362# a_4584_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X128 a_6852_n2362# a_6852_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X129 a_3828_n2362# a_3828_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X130 a_n2598_1394# a_n2598_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X131 a_n708_n2362# a_n708_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X132 a_n4866_1394# a_n4866_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X133 a_n6756_5150# a_n6756_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X134 a_1182_n2362# a_1182_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X135 a_n6000_n2362# a_n6000_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X136 a_7230_5150# a_7230_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X137 a_3450_n2362# a_3450_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X138 a_n1464_1394# a_n1464_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X139 a_4584_5150# a_4584_1930# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X140 a_n2598_n2362# a_n2598_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X141 a_n3732_1394# a_n3732_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X142 a_n4866_n2362# a_n4866_n5582# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X143 a_426_1394# a_426_n1826# 0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
C0 a_n4866_n2362# a_n4488_n2362# 0.296258f
C1 a_48_1394# a_48_1930# 0.180952f
C2 a_7230_5150# a_7608_5150# 0.296258f
C3 a_5718_1394# a_5340_1394# 0.296258f
C4 a_n2976_1930# a_n3354_1930# 0.296258f
C5 a_2316_1394# a_2694_1394# 0.296258f
C6 a_n1464_1394# a_n1842_1394# 0.296258f
C7 a_2694_n2362# a_2316_n2362# 0.296258f
C8 a_n1464_n1826# a_n1086_n1826# 0.296258f
C9 a_3828_n5582# a_3450_n5582# 0.296258f
C10 a_n5622_1394# a_n6000_1394# 0.296258f
C11 a_4206_n5582# a_4584_n5582# 0.296258f
C12 a_7230_n2362# a_6852_n2362# 0.296258f
C13 a_n2976_n2362# a_n2598_n2362# 0.296258f
C14 a_7986_1930# a_7608_1930# 0.296258f
C15 a_n7512_1394# a_n7134_1394# 0.296258f
C16 a_8742_5150# a_8364_5150# 0.296258f
C17 a_4962_5150# a_4584_5150# 0.296258f
C18 a_1182_n1826# a_1560_n1826# 0.296258f
C19 a_426_1930# a_48_1930# 0.296258f
C20 a_n7134_n1826# a_n6756_n1826# 0.296258f
C21 a_4962_n1826# a_4584_n1826# 0.296258f
C22 a_n3354_n5582# a_n2976_n5582# 0.296258f
C23 a_n2220_n2362# a_n2220_n1826# 0.180952f
C24 a_804_n2362# a_1182_n2362# 0.296258f
C25 a_48_n1826# a_n330_n1826# 0.296258f
C26 a_7230_n1826# a_6852_n1826# 0.296258f
C27 a_n2976_1394# a_n2976_1930# 0.180952f
C28 a_n1842_n5582# a_n1464_n5582# 0.296258f
C29 a_3450_n1826# a_3450_n2362# 0.180952f
C30 a_4206_n1826# a_4584_n1826# 0.296258f
C31 a_n4110_n2362# a_n4110_n1826# 0.180952f
C32 a_1182_n1826# a_1182_n2362# 0.180952f
C33 a_n7512_5150# a_n7134_5150# 0.296258f
C34 a_3828_n1826# a_3450_n1826# 0.296258f
C35 a_n6000_n5582# a_n6378_n5582# 0.296258f
C36 a_n8268_1394# a_n8646_1394# 0.296258f
C37 a_n708_n2362# a_n708_n1826# 0.180952f
C38 a_n9024_1394# a_n9024_1930# 0.180952f
C39 a_n708_1394# a_n330_1394# 0.296258f
C40 a_1938_1394# a_1938_1930# 0.180952f
C41 a_n5622_n5582# a_n5244_n5582# 0.296258f
C42 a_n7890_n1826# a_n8268_n1826# 0.296258f
C43 a_3072_n1826# a_3072_n2362# 0.180952f
C44 a_3450_5150# a_3072_5150# 0.296258f
C45 a_n2598_n5582# a_n2220_n5582# 0.296258f
C46 a_n6378_1930# a_n6756_1930# 0.296258f
C47 a_n4110_n2362# a_n4488_n2362# 0.296258f
C48 a_6096_1394# a_6474_1394# 0.296258f
C49 a_n8268_1930# a_n7890_1930# 0.296258f
C50 a_n4110_1930# a_n4488_1930# 0.296258f
C51 a_1938_1394# a_1560_1394# 0.296258f
C52 a_3450_1930# a_3828_1930# 0.296258f
C53 a_n4866_n2362# a_n4866_n1826# 0.180952f
C54 a_4206_1394# a_4206_1930# 0.180952f
C55 a_n330_1930# a_n330_1394# 0.180952f
C56 a_2694_n1826# a_2316_n1826# 0.296258f
C57 a_48_1394# a_n330_1394# 0.296258f
C58 a_n6756_n2362# a_n6756_n1826# 0.180952f
C59 a_n5622_n2362# a_n5622_n1826# 0.180952f
C60 a_n6378_n2362# a_n6000_n2362# 0.296258f
C61 a_n1842_1930# a_n2220_1930# 0.296258f
C62 a_3072_n2362# a_2694_n2362# 0.296258f
C63 a_n6000_n2362# a_n6000_n1826# 0.180952f
C64 a_n4866_1930# a_n4866_1394# 0.180952f
C65 a_n8268_5150# a_n8646_5150# 0.296258f
C66 a_5718_1394# a_6096_1394# 0.296258f
C67 a_4584_1930# a_4206_1930# 0.296258f
C68 a_n708_1394# a_n708_1930# 0.180952f
C69 a_n1842_n2362# a_n2220_n2362# 0.296258f
C70 a_48_5150# a_426_5150# 0.296258f
C71 a_4584_n2362# a_4962_n2362# 0.296258f
C72 a_n2976_n2362# a_n3354_n2362# 0.296258f
C73 a_n1842_n5582# a_n2220_n5582# 0.296258f
C74 a_5340_5150# a_5718_5150# 0.296258f
C75 a_6474_n1826# a_6852_n1826# 0.296258f
C76 a_6852_n1826# a_6852_n2362# 0.180952f
C77 a_n9024_5150# a_n8646_5150# 0.296258f
C78 a_8364_n5582# a_7986_n5582# 0.296258f
C79 a_804_n2362# a_426_n2362# 0.296258f
C80 a_n8268_1930# a_n8646_1930# 0.296258f
C81 a_4962_n5582# a_4584_n5582# 0.296258f
C82 a_n2220_n2362# a_n2598_n2362# 0.296258f
C83 a_5340_1394# a_5340_1930# 0.180952f
C84 a_n330_1930# a_n708_1930# 0.296258f
C85 a_1182_n5582# a_804_n5582# 0.296258f
C86 a_n3354_5150# a_n2976_5150# 0.296258f
C87 a_n5244_5150# a_n4866_5150# 0.296258f
C88 a_n4866_n5582# a_n5244_n5582# 0.296258f
C89 a_3828_5150# a_4206_5150# 0.296258f
C90 a_7986_1394# a_8364_1394# 0.296258f
C91 a_n2598_n5582# a_n2976_n5582# 0.296258f
C92 a_5340_1394# a_4962_1394# 0.296258f
C93 a_n1464_n2362# a_n1842_n2362# 0.296258f
C94 a_3828_1930# a_3828_1394# 0.180952f
C95 a_n1464_1394# a_n1464_1930# 0.180952f
C96 a_1938_n5582# a_2316_n5582# 0.296258f
C97 a_6474_1930# a_6474_1394# 0.180952f
C98 a_n2220_n1826# a_n2598_n1826# 0.296258f
C99 a_n7890_n5582# a_n7512_n5582# 0.296258f
C100 a_4584_1394# a_4962_1394# 0.296258f
C101 a_n8646_n2362# a_n8646_n1826# 0.180952f
C102 a_5718_n5582# a_6096_n5582# 0.296258f
C103 a_2316_1930# a_2316_1394# 0.180952f
C104 a_2694_1930# a_2694_1394# 0.180952f
C105 a_48_5150# a_n330_5150# 0.296258f
C106 a_n3354_n5582# a_n3732_n5582# 0.296258f
C107 a_4962_n5582# a_5340_n5582# 0.296258f
C108 a_7986_5150# a_7608_5150# 0.296258f
C109 a_426_1930# a_804_1930# 0.296258f
C110 a_n6378_5150# a_n6756_5150# 0.296258f
C111 a_n6000_n2362# a_n5622_n2362# 0.296258f
C112 a_804_5150# a_426_5150# 0.296258f
C113 a_n7890_n1826# a_n7512_n1826# 0.296258f
C114 a_n6378_n2362# a_n6378_n1826# 0.180952f
C115 a_n7512_n1826# a_n7512_n2362# 0.180952f
C116 a_n8268_n5582# a_n7890_n5582# 0.296258f
C117 a_n1086_n5582# a_n1464_n5582# 0.296258f
C118 a_n6000_n1826# a_n6378_n1826# 0.296258f
C119 a_n5622_n5582# a_n6000_n5582# 0.296258f
C120 a_426_n5582# a_48_n5582# 0.296258f
C121 a_n1842_1930# a_n1842_1394# 0.180952f
C122 a_n2976_n2362# a_n2976_n1826# 0.180952f
C123 a_5340_n2362# a_4962_n2362# 0.296258f
C124 a_n3732_1930# a_n3732_1394# 0.180952f
C125 a_3072_5150# a_2694_5150# 0.296258f
C126 a_426_1394# a_48_1394# 0.296258f
C127 a_n1086_n1826# a_n1086_n2362# 0.180952f
C128 a_n1086_5150# a_n1464_5150# 0.296258f
C129 a_n8646_1394# a_n8646_1930# 0.180952f
C130 a_2694_n5582# a_2316_n5582# 0.296258f
C131 a_7608_1930# a_7608_1394# 0.180952f
C132 a_4584_n2362# a_4206_n2362# 0.296258f
C133 a_n9024_n2362# a_n9024_n1826# 0.180952f
C134 a_6096_n5582# a_6474_n5582# 0.296258f
C135 a_n4488_1394# a_n4866_1394# 0.296258f
C136 a_6852_1394# a_6474_1394# 0.296258f
C137 a_7608_n1826# a_7986_n1826# 0.296258f
C138 a_n3732_n2362# a_n4110_n2362# 0.296258f
C139 a_2316_1930# a_1938_1930# 0.296258f
C140 a_n2598_n2362# a_n2598_n1826# 0.180952f
C141 a_7230_1394# a_7230_1930# 0.180952f
C142 a_6096_1394# a_6096_1930# 0.180952f
C143 a_7608_n2362# a_7986_n2362# 0.296258f
C144 a_n5244_n1826# a_n5622_n1826# 0.296258f
C145 a_7986_5150# a_8364_5150# 0.296258f
C146 a_n1086_n5582# a_n708_n5582# 0.296258f
C147 a_4962_5150# a_5340_5150# 0.296258f
C148 a_426_1394# a_426_1930# 0.180952f
C149 a_n2220_1930# a_n2598_1930# 0.296258f
C150 a_804_n2362# a_804_n1826# 0.180952f
C151 a_n8268_n2362# a_n7890_n2362# 0.296258f
C152 a_n6756_1394# a_n7134_1394# 0.296258f
C153 a_3072_n2362# a_3450_n2362# 0.296258f
C154 a_n2220_1930# a_n2220_1394# 0.180952f
C155 a_3450_n5582# a_3072_n5582# 0.296258f
C156 a_8364_n1826# a_8364_n2362# 0.180952f
C157 a_n3732_n1826# a_n4110_n1826# 0.296258f
C158 a_n8646_n2362# a_n8268_n2362# 0.296258f
C159 a_n3354_1394# a_n3732_1394# 0.296258f
C160 a_3072_1394# a_3072_1930# 0.180952f
C161 a_8742_n2362# a_8364_n2362# 0.296258f
C162 a_804_n1826# a_1182_n1826# 0.296258f
C163 a_n2598_5150# a_n2976_5150# 0.296258f
C164 a_7986_1930# a_7986_1394# 0.180952f
C165 a_n6756_1394# a_n6756_1930# 0.180952f
C166 a_n708_n2362# a_n330_n2362# 0.296258f
C167 a_n7134_n2362# a_n7512_n2362# 0.296258f
C168 a_6474_1930# a_6852_1930# 0.296258f
C169 a_n1464_n2362# a_n1464_n1826# 0.180952f
C170 a_n5244_1394# a_n5244_1930# 0.180952f
C171 a_4584_1930# a_4962_1930# 0.296258f
C172 a_3828_5150# a_3450_5150# 0.296258f
C173 a_n3732_1930# a_n3354_1930# 0.296258f
C174 a_804_1930# a_1182_1930# 0.296258f
C175 a_n1086_n1826# a_n708_n1826# 0.296258f
C176 a_8364_1930# a_8364_1394# 0.180952f
C177 a_n4488_n5582# a_n4866_n5582# 0.296258f
C178 a_5718_n2362# a_5340_n2362# 0.296258f
C179 a_1182_1394# a_1182_1930# 0.180952f
C180 a_2316_1930# a_2694_1930# 0.296258f
C181 a_6096_5150# a_5718_5150# 0.296258f
C182 a_6474_5150# a_6096_5150# 0.296258f
C183 a_3450_1930# a_3072_1930# 0.296258f
C184 a_6474_1930# a_6096_1930# 0.296258f
C185 a_7986_n2362# a_8364_n2362# 0.296258f
C186 a_426_n5582# a_804_n5582# 0.296258f
C187 a_5718_1930# a_5718_1394# 0.180952f
C188 a_1560_1930# a_1182_1930# 0.296258f
C189 a_4584_5150# a_4206_5150# 0.296258f
C190 a_n4110_1394# a_n3732_1394# 0.296258f
C191 a_n8268_1394# a_n7890_1394# 0.296258f
C192 a_1938_n1826# a_2316_n1826# 0.296258f
C193 a_3828_1930# a_4206_1930# 0.296258f
C194 a_n330_n1826# a_n708_n1826# 0.296258f
C195 a_2316_n2362# a_2316_n1826# 0.180952f
C196 a_n7134_n5582# a_n6756_n5582# 0.296258f
C197 a_n3354_1394# a_n3354_1930# 0.180952f
C198 a_n3354_5150# a_n3732_5150# 0.296258f
C199 a_426_n2362# a_426_n1826# 0.180952f
C200 a_n1842_1930# a_n1464_1930# 0.296258f
C201 a_8742_1394# a_8364_1394# 0.296258f
C202 a_n1842_5150# a_n2220_5150# 0.296258f
C203 a_n6000_1930# a_n5622_1930# 0.296258f
C204 a_n5244_n2362# a_n5622_n2362# 0.296258f
C205 a_5340_n1826# a_5340_n2362# 0.180952f
C206 a_n330_n5582# a_n708_n5582# 0.296258f
C207 a_4962_n1826# a_4962_n2362# 0.180952f
C208 a_6852_1394# a_6852_1930# 0.180952f
C209 a_n3354_n1826# a_n3732_n1826# 0.296258f
C210 a_n1842_1394# a_n2220_1394# 0.296258f
C211 a_n2976_1394# a_n3354_1394# 0.296258f
C212 a_n5622_1930# a_n5244_1930# 0.296258f
C213 a_48_n2362# a_n330_n2362# 0.296258f
C214 a_n4866_1930# a_n4488_1930# 0.296258f
C215 a_6852_5150# a_7230_5150# 0.296258f
C216 a_8364_1930# a_8742_1930# 0.296258f
C217 a_n9024_n5582# a_n8646_n5582# 0.296258f
C218 a_n8646_n1826# a_n8268_n1826# 0.296258f
C219 a_n3354_n1826# a_n3354_n2362# 0.180952f
C220 a_426_n2362# a_48_n2362# 0.296258f
C221 a_1560_1930# a_1938_1930# 0.296258f
C222 a_1560_1394# a_1182_1394# 0.296258f
C223 a_n6378_1394# a_n6000_1394# 0.296258f
C224 a_3072_n1826# a_2694_n1826# 0.296258f
C225 a_n7512_1930# a_n7890_1930# 0.296258f
C226 a_1560_1394# a_1560_1930# 0.180952f
C227 a_n6378_1930# a_n6378_1394# 0.180952f
C228 a_n7134_n1826# a_n7512_n1826# 0.296258f
C229 a_3828_n2362# a_4206_n2362# 0.296258f
C230 a_n1086_1394# a_n1086_1930# 0.180952f
C231 a_n2976_n1826# a_n2598_n1826# 0.296258f
C232 a_8742_1930# a_8742_1394# 0.180952f
C233 a_7986_1930# a_8364_1930# 0.296258f
C234 a_n7134_n5582# a_n7512_n5582# 0.296258f
C235 a_2694_n2362# a_2694_n1826# 0.180952f
C236 a_7230_n5582# a_6852_n5582# 0.296258f
C237 a_2694_1394# a_3072_1394# 0.296258f
C238 a_n8646_1394# a_n9024_1394# 0.296258f
C239 a_n4110_1394# a_n4488_1394# 0.296258f
C240 a_n2598_1394# a_n2598_1930# 0.180952f
C241 a_n2598_1394# a_n2220_1394# 0.296258f
C242 a_4584_n2362# a_4584_n1826# 0.180952f
C243 a_n3732_n2362# a_n3732_n1826# 0.180952f
C244 a_5718_1930# a_5340_1930# 0.296258f
C245 a_n7890_1394# a_n7890_1930# 0.180952f
C246 a_n1842_n1826# a_n2220_n1826# 0.296258f
C247 a_n6000_1930# a_n6000_1394# 0.180952f
C248 a_7608_1394# a_7986_1394# 0.296258f
C249 a_7608_n5582# a_7230_n5582# 0.296258f
C250 a_n4110_n5582# a_n4488_n5582# 0.296258f
C251 a_n6756_n2362# a_n6378_n2362# 0.296258f
C252 a_1182_n5582# a_1560_n5582# 0.296258f
C253 a_804_n1826# a_426_n1826# 0.296258f
C254 a_n6000_1930# a_n6378_1930# 0.296258f
C255 a_n3732_n2362# a_n3354_n2362# 0.296258f
C256 a_n5622_1394# a_n5244_1394# 0.296258f
C257 a_48_n1826# a_426_n1826# 0.296258f
C258 a_5718_1930# a_6096_1930# 0.296258f
C259 a_8742_n5582# a_8364_n5582# 0.296258f
C260 a_n330_n5582# a_48_n5582# 0.296258f
C261 a_n6756_n1826# a_n6378_n1826# 0.296258f
C262 a_n4866_1394# a_n5244_1394# 0.296258f
C263 a_n1464_n2362# a_n1086_n2362# 0.296258f
C264 a_n7890_n1826# a_n7890_n2362# 0.180952f
C265 a_n7512_n2362# a_n7890_n2362# 0.296258f
C266 a_n6756_5150# a_n7134_5150# 0.296258f
C267 a_4206_n5582# a_3828_n5582# 0.296258f
C268 a_1182_5150# a_1560_5150# 0.296258f
C269 a_1560_n2362# a_1560_n1826# 0.180952f
C270 a_n3354_n1826# a_n2976_n1826# 0.296258f
C271 a_4206_n1826# a_4206_n2362# 0.180952f
C272 a_n7512_1930# a_n7134_1930# 0.296258f
C273 a_n8268_5150# a_n7890_5150# 0.296258f
C274 a_4584_1394# a_4206_1394# 0.296258f
C275 a_n8268_n1826# a_n8268_n2362# 0.180952f
C276 a_6096_n2362# a_6474_n2362# 0.296258f
C277 a_6096_n1826# a_5718_n1826# 0.296258f
C278 a_n7134_n1826# a_n7134_n2362# 0.180952f
C279 a_1938_5150# a_1560_5150# 0.296258f
C280 a_n5244_n2362# a_n5244_n1826# 0.180952f
C281 a_n2976_1394# a_n2598_1394# 0.296258f
C282 a_5340_n1826# a_4962_n1826# 0.296258f
C283 a_1560_n2362# a_1182_n2362# 0.296258f
C284 a_4584_1394# a_4584_1930# 0.180952f
C285 a_n8646_1930# a_n9024_1930# 0.296258f
C286 a_n2220_5150# a_n2598_5150# 0.296258f
C287 a_n4488_1394# a_n4488_1930# 0.180952f
C288 a_5718_n5582# a_5340_n5582# 0.296258f
C289 a_n8646_n2362# a_n9024_n2362# 0.296258f
C290 a_3072_n1826# a_3450_n1826# 0.296258f
C291 a_1560_n2362# a_1938_n2362# 0.296258f
C292 a_n8646_n1826# a_n9024_n1826# 0.296258f
C293 a_n1842_n2362# a_n1842_n1826# 0.180952f
C294 a_48_n1826# a_48_n2362# 0.180952f
C295 a_n4488_n1826# a_n4110_n1826# 0.296258f
C296 a_7608_n1826# a_7608_n2362# 0.180952f
C297 a_n4110_n5582# a_n3732_n5582# 0.296258f
C298 a_6852_n5582# a_6474_n5582# 0.296258f
C299 a_5718_n2362# a_5718_n1826# 0.180952f
C300 a_3072_1394# a_3450_1394# 0.296258f
C301 a_7608_n5582# a_7986_n5582# 0.296258f
C302 a_7608_1930# a_7230_1930# 0.296258f
C303 a_n330_n1826# a_n330_n2362# 0.180952f
C304 a_8364_n1826# a_7986_n1826# 0.296258f
C305 a_n7512_1930# a_n7512_1394# 0.180952f
C306 a_n6000_5150# a_n5622_5150# 0.296258f
C307 a_n4110_1930# a_n3732_1930# 0.296258f
C308 a_n4488_n2362# a_n4488_n1826# 0.180952f
C309 a_n4866_1930# a_n5244_1930# 0.296258f
C310 a_n6756_n2362# a_n7134_n2362# 0.296258f
C311 a_7230_n1826# a_7608_n1826# 0.296258f
C312 a_4206_1394# a_3828_1394# 0.296258f
C313 a_3828_n2362# a_3450_n2362# 0.296258f
C314 a_n4488_5150# a_n4110_5150# 0.296258f
C315 a_n5622_1930# a_n5622_1394# 0.180952f
C316 a_6474_n2362# a_6474_n1826# 0.180952f
C317 a_6474_n2362# a_6852_n2362# 0.296258f
C318 a_1938_n5582# a_1560_n5582# 0.296258f
C319 a_3828_n1826# a_3828_n2362# 0.180952f
C320 a_2316_5150# a_2694_5150# 0.296258f
C321 a_7608_n2362# a_7230_n2362# 0.296258f
C322 a_4962_1930# a_5340_1930# 0.296258f
C323 a_n1086_1930# a_n708_1930# 0.296258f
C324 a_7608_1394# a_7230_1394# 0.296258f
C325 a_n1464_1394# a_n1086_1394# 0.296258f
C326 a_1938_n1826# a_1560_n1826# 0.296258f
C327 a_n3732_5150# a_n4110_5150# 0.296258f
C328 a_4962_1930# a_4962_1394# 0.180952f
C329 a_6096_n2362# a_6096_n1826# 0.180952f
C330 a_n7512_1394# a_n7890_1394# 0.296258f
C331 a_5340_n1826# a_5718_n1826# 0.296258f
C332 a_n4866_n2362# a_n5244_n2362# 0.296258f
C333 a_n4488_5150# a_n4866_5150# 0.296258f
C334 a_804_1930# a_804_1394# 0.180952f
C335 a_3450_1930# a_3450_1394# 0.180952f
C336 a_n1086_1394# a_n708_1394# 0.296258f
C337 a_n1086_5150# a_n708_5150# 0.296258f
C338 a_804_1394# a_1182_1394# 0.296258f
C339 a_8364_n1826# a_8742_n1826# 0.296258f
C340 a_2694_n5582# a_3072_n5582# 0.296258f
C341 a_n8268_1394# a_n8268_1930# 0.180952f
C342 a_8742_n2362# a_8742_n1826# 0.180952f
C343 a_7230_n1826# a_7230_n2362# 0.180952f
C344 a_7986_n2362# a_7986_n1826# 0.180952f
C345 a_7230_1930# a_6852_1930# 0.296258f
C346 a_6852_5150# a_6474_5150# 0.296258f
C347 a_n6756_1394# a_n6378_1394# 0.296258f
C348 a_1938_n1826# a_1938_n2362# 0.180952f
C349 a_n708_5150# a_n330_5150# 0.296258f
C350 a_n6378_n5582# a_n6756_n5582# 0.296258f
C351 a_n6378_5150# a_n6000_5150# 0.296258f
C352 a_2316_n2362# a_1938_n2362# 0.296258f
C353 a_804_5150# a_1182_5150# 0.296258f
C354 a_n8268_n5582# a_n8646_n5582# 0.296258f
C355 a_6096_n2362# a_5718_n2362# 0.296258f
C356 a_n1842_5150# a_n1464_5150# 0.296258f
C357 a_n7134_1394# a_n7134_1930# 0.180952f
C358 a_2316_1394# a_1938_1394# 0.296258f
C359 a_n4866_n1826# a_n4488_n1826# 0.296258f
C360 a_n2976_1930# a_n2598_1930# 0.296258f
C361 a_n708_n2362# a_n1086_n2362# 0.296258f
C362 a_n7512_5150# a_n7890_5150# 0.296258f
C363 a_4206_n1826# a_3828_n1826# 0.296258f
C364 a_n1086_1930# a_n1464_1930# 0.296258f
C365 a_n7134_1930# a_n6756_1930# 0.296258f
C366 a_n6000_n1826# a_n5622_n1826# 0.296258f
C367 a_7230_1394# a_6852_1394# 0.296258f
C368 a_n5244_5150# a_n5622_5150# 0.296258f
C369 a_426_1394# a_804_1394# 0.296258f
C370 a_n4866_n1826# a_n5244_n1826# 0.296258f
C371 a_2694_1930# a_3072_1930# 0.296258f
C372 a_3828_1394# a_3450_1394# 0.296258f
C373 a_n1464_n1826# a_n1842_n1826# 0.296258f
C374 a_6096_n1826# a_6474_n1826# 0.296258f
C375 a_n4110_1930# a_n4110_1394# 0.180952f
C376 a_1938_5150# a_2316_5150# 0.296258f
C377 a_n330_1930# a_48_1930# 0.296258f
C378 a_8742_n5582# 0 0.626416f
C379 a_8742_n2362# 0 0.494677f
C380 a_8364_n5582# 0 0.417886f
C381 a_8364_n2362# 0 0.286147f
C382 a_7986_n5582# 0 0.417886f
C383 a_7986_n2362# 0 0.286147f
C384 a_7608_n5582# 0 0.417886f
C385 a_7608_n2362# 0 0.286147f
C386 a_7230_n5582# 0 0.417886f
C387 a_7230_n2362# 0 0.286147f
C388 a_6852_n5582# 0 0.417886f
C389 a_6852_n2362# 0 0.286147f
C390 a_6474_n5582# 0 0.417886f
C391 a_6474_n2362# 0 0.286147f
C392 a_6096_n5582# 0 0.417886f
C393 a_6096_n2362# 0 0.286147f
C394 a_5718_n5582# 0 0.417886f
C395 a_5718_n2362# 0 0.286147f
C396 a_5340_n5582# 0 0.417886f
C397 a_5340_n2362# 0 0.286147f
C398 a_4962_n5582# 0 0.417886f
C399 a_4962_n2362# 0 0.286147f
C400 a_4584_n5582# 0 0.417886f
C401 a_4584_n2362# 0 0.286147f
C402 a_4206_n5582# 0 0.417886f
C403 a_4206_n2362# 0 0.286147f
C404 a_3828_n5582# 0 0.417886f
C405 a_3828_n2362# 0 0.286147f
C406 a_3450_n5582# 0 0.417886f
C407 a_3450_n2362# 0 0.286147f
C408 a_3072_n5582# 0 0.417886f
C409 a_3072_n2362# 0 0.286147f
C410 a_2694_n5582# 0 0.417886f
C411 a_2694_n2362# 0 0.286147f
C412 a_2316_n5582# 0 0.417886f
C413 a_2316_n2362# 0 0.286147f
C414 a_1938_n5582# 0 0.417886f
C415 a_1938_n2362# 0 0.286147f
C416 a_1560_n5582# 0 0.417886f
C417 a_1560_n2362# 0 0.286147f
C418 a_1182_n5582# 0 0.417886f
C419 a_1182_n2362# 0 0.286147f
C420 a_804_n5582# 0 0.417886f
C421 a_804_n2362# 0 0.286147f
C422 a_426_n5582# 0 0.417886f
C423 a_426_n2362# 0 0.286147f
C424 a_48_n5582# 0 0.417886f
C425 a_48_n2362# 0 0.286147f
C426 a_n330_n5582# 0 0.417886f
C427 a_n330_n2362# 0 0.286147f
C428 a_n708_n5582# 0 0.417886f
C429 a_n708_n2362# 0 0.286147f
C430 a_n1086_n5582# 0 0.417886f
C431 a_n1086_n2362# 0 0.286147f
C432 a_n1464_n5582# 0 0.417886f
C433 a_n1464_n2362# 0 0.286147f
C434 a_n1842_n5582# 0 0.417886f
C435 a_n1842_n2362# 0 0.286147f
C436 a_n2220_n5582# 0 0.417886f
C437 a_n2220_n2362# 0 0.286147f
C438 a_n2598_n5582# 0 0.417886f
C439 a_n2598_n2362# 0 0.286147f
C440 a_n2976_n5582# 0 0.417886f
C441 a_n2976_n2362# 0 0.286147f
C442 a_n3354_n5582# 0 0.417886f
C443 a_n3354_n2362# 0 0.286147f
C444 a_n3732_n5582# 0 0.417886f
C445 a_n3732_n2362# 0 0.286147f
C446 a_n4110_n5582# 0 0.417886f
C447 a_n4110_n2362# 0 0.286147f
C448 a_n4488_n5582# 0 0.417886f
C449 a_n4488_n2362# 0 0.286147f
C450 a_n4866_n5582# 0 0.417886f
C451 a_n4866_n2362# 0 0.286147f
C452 a_n5244_n5582# 0 0.417886f
C453 a_n5244_n2362# 0 0.286147f
C454 a_n5622_n5582# 0 0.417886f
C455 a_n5622_n2362# 0 0.286147f
C456 a_n6000_n5582# 0 0.417886f
C457 a_n6000_n2362# 0 0.286147f
C458 a_n6378_n5582# 0 0.417886f
C459 a_n6378_n2362# 0 0.286147f
C460 a_n6756_n5582# 0 0.417886f
C461 a_n6756_n2362# 0 0.286147f
C462 a_n7134_n5582# 0 0.417886f
C463 a_n7134_n2362# 0 0.286147f
C464 a_n7512_n5582# 0 0.417886f
C465 a_n7512_n2362# 0 0.286147f
C466 a_n7890_n5582# 0 0.417886f
C467 a_n7890_n2362# 0 0.286147f
C468 a_n8268_n5582# 0 0.417886f
C469 a_n8268_n2362# 0 0.286147f
C470 a_n8646_n5582# 0 0.417886f
C471 a_n8646_n2362# 0 0.286147f
C472 a_n9024_n5582# 0 0.626416f
C473 a_n9024_n2362# 0 0.494677f
C474 a_8742_n1826# 0 0.494677f
C475 a_8742_1394# 0 0.494677f
C476 a_8364_n1826# 0 0.286147f
C477 a_8364_1394# 0 0.286147f
C478 a_7986_n1826# 0 0.286147f
C479 a_7986_1394# 0 0.286147f
C480 a_7608_n1826# 0 0.286147f
C481 a_7608_1394# 0 0.286147f
C482 a_7230_n1826# 0 0.286147f
C483 a_7230_1394# 0 0.286147f
C484 a_6852_n1826# 0 0.286147f
C485 a_6852_1394# 0 0.286147f
C486 a_6474_n1826# 0 0.286147f
C487 a_6474_1394# 0 0.286147f
C488 a_6096_n1826# 0 0.286147f
C489 a_6096_1394# 0 0.286147f
C490 a_5718_n1826# 0 0.286147f
C491 a_5718_1394# 0 0.286147f
C492 a_5340_n1826# 0 0.286147f
C493 a_5340_1394# 0 0.286147f
C494 a_4962_n1826# 0 0.286147f
C495 a_4962_1394# 0 0.286147f
C496 a_4584_n1826# 0 0.286147f
C497 a_4584_1394# 0 0.286147f
C498 a_4206_n1826# 0 0.286147f
C499 a_4206_1394# 0 0.286147f
C500 a_3828_n1826# 0 0.286147f
C501 a_3828_1394# 0 0.286147f
C502 a_3450_n1826# 0 0.286147f
C503 a_3450_1394# 0 0.286147f
C504 a_3072_n1826# 0 0.286147f
C505 a_3072_1394# 0 0.286147f
C506 a_2694_n1826# 0 0.286147f
C507 a_2694_1394# 0 0.286147f
C508 a_2316_n1826# 0 0.286147f
C509 a_2316_1394# 0 0.286147f
C510 a_1938_n1826# 0 0.286147f
C511 a_1938_1394# 0 0.286147f
C512 a_1560_n1826# 0 0.286147f
C513 a_1560_1394# 0 0.286147f
C514 a_1182_n1826# 0 0.286147f
C515 a_1182_1394# 0 0.286147f
C516 a_804_n1826# 0 0.286147f
C517 a_804_1394# 0 0.286147f
C518 a_426_n1826# 0 0.286147f
C519 a_426_1394# 0 0.286147f
C520 a_48_n1826# 0 0.286147f
C521 a_48_1394# 0 0.286147f
C522 a_n330_n1826# 0 0.286147f
C523 a_n330_1394# 0 0.286147f
C524 a_n708_n1826# 0 0.286147f
C525 a_n708_1394# 0 0.286147f
C526 a_n1086_n1826# 0 0.286147f
C527 a_n1086_1394# 0 0.286147f
C528 a_n1464_n1826# 0 0.286147f
C529 a_n1464_1394# 0 0.286147f
C530 a_n1842_n1826# 0 0.286147f
C531 a_n1842_1394# 0 0.286147f
C532 a_n2220_n1826# 0 0.286147f
C533 a_n2220_1394# 0 0.286147f
C534 a_n2598_n1826# 0 0.286147f
C535 a_n2598_1394# 0 0.286147f
C536 a_n2976_n1826# 0 0.286147f
C537 a_n2976_1394# 0 0.286147f
C538 a_n3354_n1826# 0 0.286147f
C539 a_n3354_1394# 0 0.286147f
C540 a_n3732_n1826# 0 0.286147f
C541 a_n3732_1394# 0 0.286147f
C542 a_n4110_n1826# 0 0.286147f
C543 a_n4110_1394# 0 0.286147f
C544 a_n4488_n1826# 0 0.286147f
C545 a_n4488_1394# 0 0.286147f
C546 a_n4866_n1826# 0 0.286147f
C547 a_n4866_1394# 0 0.286147f
C548 a_n5244_n1826# 0 0.286147f
C549 a_n5244_1394# 0 0.286147f
C550 a_n5622_n1826# 0 0.286147f
C551 a_n5622_1394# 0 0.286147f
C552 a_n6000_n1826# 0 0.286147f
C553 a_n6000_1394# 0 0.286147f
C554 a_n6378_n1826# 0 0.286147f
C555 a_n6378_1394# 0 0.286147f
C556 a_n6756_n1826# 0 0.286147f
C557 a_n6756_1394# 0 0.286147f
C558 a_n7134_n1826# 0 0.286147f
C559 a_n7134_1394# 0 0.286147f
C560 a_n7512_n1826# 0 0.286147f
C561 a_n7512_1394# 0 0.286147f
C562 a_n7890_n1826# 0 0.286147f
C563 a_n7890_1394# 0 0.286147f
C564 a_n8268_n1826# 0 0.286147f
C565 a_n8268_1394# 0 0.286147f
C566 a_n8646_n1826# 0 0.286147f
C567 a_n8646_1394# 0 0.286147f
C568 a_n9024_n1826# 0 0.494677f
C569 a_n9024_1394# 0 0.494677f
C570 a_8742_1930# 0 0.494677f
C571 a_8742_5150# 0 0.626416f
C572 a_8364_1930# 0 0.286147f
C573 a_8364_5150# 0 0.417886f
C574 a_7986_1930# 0 0.286147f
C575 a_7986_5150# 0 0.417886f
C576 a_7608_1930# 0 0.286147f
C577 a_7608_5150# 0 0.417886f
C578 a_7230_1930# 0 0.286147f
C579 a_7230_5150# 0 0.417886f
C580 a_6852_1930# 0 0.286147f
C581 a_6852_5150# 0 0.417886f
C582 a_6474_1930# 0 0.286147f
C583 a_6474_5150# 0 0.417886f
C584 a_6096_1930# 0 0.286147f
C585 a_6096_5150# 0 0.417886f
C586 a_5718_1930# 0 0.286147f
C587 a_5718_5150# 0 0.417886f
C588 a_5340_1930# 0 0.286147f
C589 a_5340_5150# 0 0.417886f
C590 a_4962_1930# 0 0.286147f
C591 a_4962_5150# 0 0.417886f
C592 a_4584_1930# 0 0.286147f
C593 a_4584_5150# 0 0.417886f
C594 a_4206_1930# 0 0.286147f
C595 a_4206_5150# 0 0.417886f
C596 a_3828_1930# 0 0.286147f
C597 a_3828_5150# 0 0.417886f
C598 a_3450_1930# 0 0.286147f
C599 a_3450_5150# 0 0.417886f
C600 a_3072_1930# 0 0.286147f
C601 a_3072_5150# 0 0.417886f
C602 a_2694_1930# 0 0.286147f
C603 a_2694_5150# 0 0.417886f
C604 a_2316_1930# 0 0.286147f
C605 a_2316_5150# 0 0.417886f
C606 a_1938_1930# 0 0.286147f
C607 a_1938_5150# 0 0.417886f
C608 a_1560_1930# 0 0.286147f
C609 a_1560_5150# 0 0.417886f
C610 a_1182_1930# 0 0.286147f
C611 a_1182_5150# 0 0.417886f
C612 a_804_1930# 0 0.286147f
C613 a_804_5150# 0 0.417886f
C614 a_426_1930# 0 0.286147f
C615 a_426_5150# 0 0.417886f
C616 a_48_1930# 0 0.286147f
C617 a_48_5150# 0 0.417886f
C618 a_n330_1930# 0 0.286147f
C619 a_n330_5150# 0 0.417886f
C620 a_n708_1930# 0 0.286147f
C621 a_n708_5150# 0 0.417886f
C622 a_n1086_1930# 0 0.286147f
C623 a_n1086_5150# 0 0.417886f
C624 a_n1464_1930# 0 0.286147f
C625 a_n1464_5150# 0 0.417886f
C626 a_n1842_1930# 0 0.286147f
C627 a_n1842_5150# 0 0.417886f
C628 a_n2220_1930# 0 0.286147f
C629 a_n2220_5150# 0 0.417886f
C630 a_n2598_1930# 0 0.286147f
C631 a_n2598_5150# 0 0.417886f
C632 a_n2976_1930# 0 0.286147f
C633 a_n2976_5150# 0 0.417886f
C634 a_n3354_1930# 0 0.286147f
C635 a_n3354_5150# 0 0.417886f
C636 a_n3732_1930# 0 0.286147f
C637 a_n3732_5150# 0 0.417886f
C638 a_n4110_1930# 0 0.286147f
C639 a_n4110_5150# 0 0.417886f
C640 a_n4488_1930# 0 0.286147f
C641 a_n4488_5150# 0 0.417886f
C642 a_n4866_1930# 0 0.286147f
C643 a_n4866_5150# 0 0.417886f
C644 a_n5244_1930# 0 0.286147f
C645 a_n5244_5150# 0 0.417886f
C646 a_n5622_1930# 0 0.286147f
C647 a_n5622_5150# 0 0.417886f
C648 a_n6000_1930# 0 0.286147f
C649 a_n6000_5150# 0 0.417886f
C650 a_n6378_1930# 0 0.286147f
C651 a_n6378_5150# 0 0.417886f
C652 a_n6756_1930# 0 0.286147f
C653 a_n6756_5150# 0 0.417886f
C654 a_n7134_1930# 0 0.286147f
C655 a_n7134_5150# 0 0.417886f
C656 a_n7512_1930# 0 0.286147f
C657 a_n7512_5150# 0 0.417886f
C658 a_n7890_1930# 0 0.286147f
C659 a_n7890_5150# 0 0.417886f
C660 a_n8268_1930# 0 0.286147f
C661 a_n8268_5150# 0 0.417886f
C662 a_n8646_1930# 0 0.286147f
C663 a_n8646_5150# 0 0.417886f
C664 a_n9024_1930# 0 0.494677f
C665 a_n9024_5150# 0 0.626416f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8 a_300_n300# a_n492_n522# a_n358_n300#
+ a_n300_n388#
X0 a_300_n300# a_n300_n388# a_n358_n300# a_n492_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=3
C0 a_n358_n300# a_300_n300# 0.064341f
C1 a_n358_n300# a_n300_n388# 0.113258f
C2 a_300_n300# a_n300_n388# 0.113258f
C3 a_300_n300# a_n492_n522# 0.381938f
C4 a_n358_n300# a_n492_n522# 0.381938f
C5 a_n300_n388# a_n492_n522# 1.81083f
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_F6RBXN a_n147_n172# a_n45_n70#
X0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
C0 a_n45_n70# a_n147_n172# 0.218219f
.ends

.subckt voltage_divider out_0000 out_0001 out_0010 out_0011 out_0101 out_0110 out_0111
+ out_1001 out_1010 out_1011 out_1101 out_1111 ena m1_7155_3601# m1_10901_8137# m1_7155_14563#
+ m1_7691_16075# m1_3399_9649# m1_10911_2089# m1_7155_3223# m1_3399_12673# m1_10911_15697#
+ m1_3399_3979# m1_7155_5491# m1_3399_7381# m1_7155_9271# m1_10911_13429# m1_7155_12295#
+ m1_7691_14563# m1_3399_16453# m1_7155_7759# m1_3935_10405# m1_179_3979# 51 m1_7155_10027#
+ m1_3399_199# m1_3399_3601# m1_179_13051# m1_3935_14185# m1_179_199# m1_7691_9271#
+ m1_7691_12295# m1_7155_10783# m1_3935_4357# m1_7691_10027# m1_7155_7003# m1_3399_15697#
+ m1_3935_8137# m1_3399_955# m1_7691_10783# m1_179_12295# m1_7155_16831# m1_179_955#
+ m1_7691_7003# m1_179_6247# m1_7155_955# m1_3399_2467# m1_179_16075# m1_3935_8893#
+ m1_3935_11917# m1_179_2467# m1_3935_5113# m1_7155_2845# m1_10911_16453# m1_3399_13429#
+ m1_7155_13051# m1_10911_1333# m1_179_16831# m1_179_10027# m1_7155_4735# m1_3399_17209#
+ m1_10911_14185# m1_179_7003# m1_3399_3223# m1_3399_6625# m1_3935_9649# m1_10911_11917#
+ m1_7691_13051# m1_179_3223# m1_3935_12673# m1_3399_2845# out_1100 m1_10911_12673#
+ m1_3935_7381# m1_3935_16453# avdd m1_7155_577# m1_7155_17209# m1_3399_5869# m1_179_10783#
+ m1_7155_199# m1_3399_11161# m1_3399_14941# m1_3399_2089# m1_7155_2467# m1_179_14563#
+ m1_7155_8515# m1_7155_15319# m1_3935_15697# m1_179_5491# m1_3399_1711# m1_7155_2089#
+ m1_179_1711# out_0100 m1_7691_15319# m1_3399_10405# m1_179_13807# m1_7155_3979#
+ m1_7155_13807# m1_3399_14185# m1_7155_6247# m1_10911_2845# m1_7155_11539# m1_179_9271#
+ m1_3399_4357# m1_3935_13429# out_1110 m1_7691_13807# m1_179_7759# m1_3399_577# m1_3399_8137#
+ out_1000 m1_3935_6625# m1_3399_8893# m1_179_11539# m1_3399_11917# m1_3399_5113#
+ m1_179_15319# m1_10911_577# m1_7155_1711# m1_7155_16075# m1_3399_1333# m1_3935_5869#
+ m1_10911_14941# m1_10901_199# m1_7155_1333# m1_179_4735# m1_179_8515# m1_3935_11161#
+ m1_3935_14941# avss
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_0 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_2 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_H3F4MM_0 m1_3399_9649# m1_7155_3979# m1_7155_16831#
+ m1_7155_2467# m1_179_955# m1_10911_577# m1_179_16831# m1_179_13051# m1_179_6247#
+ m1_179_10027# m1_3399_17209# m1_3399_2467# m1_7155_3979# m1_7155_2089# m1_179_16831#
+ m1_179_2467# m1_7155_6247# m1_10911_2845# out_1110 m1_3935_5113# m1_7155_16831#
+ m1_3935_12673# out_0011 m1_10911_15697# m1_10911_16453# m1_7155_5491# out_1110 m1_3399_1333#
+ m1_3935_4357# m1_3935_9649# m1_3935_16453# m1_3935_12673# m1_7155_13051# m1_3399_6625#
+ out_1101 out_0010 out_1000 m1_3399_8893# m1_3399_10405# m1_10911_14185# m1_179_7003#
+ m1_10911_14185# m1_179_8515# m1_179_10783# m1_3399_3223# out_1010 m1_3399_6625#
+ m1_3399_14185# m1_10911_11917# m1_3399_11161# avss m1_3399_14941# m1_7155_10783#
+ m1_7691_13051# out_0111 m1_179_3223# m1_179_6247# m1_179_14563# m1_179_10783# m1_3935_15697#
+ m1_3399_2845# m1_179_14563# m1_3399_3979# m1_3935_11917# m1_10911_11917# m1_10911_12673#
+ m1_3935_7381# m1_10911_577# m1_179_2467# out_0010 m1_7155_1711# avss m1_7691_10783#
+ m1_3399_199# m1_3935_15697# m1_3399_3601# m1_7155_17209# m1_3399_13429# m1_3399_5869#
+ m1_3399_10405# m1_10901_199# out_0001 m1_7155_1333# out_0001 m1_7155_14563# avss
+ m1_179_13807# m1_179_5491# m1_10911_2089# m1_7155_3601# m1_7155_1711# m1_179_10027#
+ avss avss m1_3399_2089# m1_3399_14185# m1_3399_5113# m1_7155_8515# m1_7155_15319#
+ m1_7155_7759# m1_7155_17209# avss m1_10911_2089# m1_179_1711# m1_7155_3223# m1_179_13807#
+ m1_7155_1333# m1_7155_8515# m1_3399_955# m1_179_5491# m1_7691_14563# m1_3399_1711#
+ m1_3935_16453# out_1101 m1_3399_8893# m1_3935_13429# m1_10911_16453# m1_7155_5491#
+ m1_3935_5869# m1_7155_15319# m1_7155_3601# avss m1_3935_9649# m1_3399_8137# m1_179_1711#
+ m1_7155_7759# m1_179_9271# m1_7155_13051# out_0100 m1_7691_15319# out_0101 m1_3399_17209#
+ out_1111 m1_7155_4735# m1_3399_2467# m1_7155_3223# out_0100 m1_179_7759# m1_3399_11161#
+ out_1001 m1_7155_7003# m1_7155_13807# out_1010 m1_7691_15319# m1_179_11539# m1_7155_11539#
+ out_0101 m1_7691_13051# m1_3399_14941# out_1001 m1_3399_4357# m1_7155_7003# out_1100
+ m1_3399_11917# m1_3399_7381# m1_10911_12673# m1_179_15319# m1_7691_7003# m1_7691_13807#
+ m1_179_3979# m1_179_11539# m1_3935_6625# m1_179_7759# m1_3399_577# m1_3935_8893#
+ m1_3935_10405# 51 m1_3399_8137# m1_7691_7003# m1_179_199# m1_3399_3223# avss m1_3935_6625#
+ out_0000 m1_3935_14185# m1_7155_955# m1_179_8515# m1_3935_11161# m1_3935_14941#
+ m1_3399_2845# m1_3399_5113# m1_10911_1333# m1_3399_12673# m1_7155_2845# m1_7155_955#
+ m1_179_4735# avdd m1_7155_9271# m1_7155_16075# m1_179_12295# m1_7155_16075# m1_3399_1333#
+ m1_10911_1333# m1_3399_4357# m1_3399_9649# m1_3399_16453# m1_3935_13429# m1_3935_5869#
+ m1_3399_12673# m1_3935_10405# m1_10911_14941# m1_179_955# out_1111 m1_7155_4735#
+ avss m1_7155_9271# m1_7155_2845# m1_179_4735# m1_179_9271# m1_179_16075# m1_179_13051#
+ avss m1_3399_2089# m1_3935_14185# m1_3935_5113# m1_10911_14941# m1_10901_8137# m1_10901_8137#
+ m1_7155_13807# m1_7691_9271# m1_7155_14563# m1_7691_16075# m1_7691_16075# m1_10911_2845#
+ out_0011 m1_7155_11539# m1_3399_1711# out_1011 m1_10911_15697# m1_7155_6247# out_1100
+ m1_7691_9271# m1_3935_8893# m1_3399_15697# m1_3399_3979# m1_3399_11917# m1_3399_7381#
+ out_0110 m1_10911_13429# m1_3935_8137# m1_7155_12295# m1_7691_13807# m1_7155_12295#
+ m1_7691_14563# out_1011 m1_179_15319# m1_179_3979# m1_179_12295# m1_179_7003# m1_7155_577#
+ m1_7155_10027# m1_3399_199# 51 m1_3399_15697# m1_3399_3601# out_0110 m1_10911_13429#
+ out_1000 m1_3935_11161# m1_179_199# m1_179_16075# out_0000 m1_7155_199# m1_179_3223#
+ m1_7155_10027# m1_7155_10783# m1_7691_12295# m1_7691_12295# avss out_0111 m1_3935_14941#
+ m1_3935_4357# m1_3935_11917# m1_7155_2467# m1_7155_577# m1_3935_7381# m1_7691_10027#
+ avss m1_3399_577# m1_3399_955# m1_7155_2089# m1_7155_199# m1_7691_10027# m1_7691_10783#
+ m1_3399_16453# avss m1_3399_13429# m1_3399_5869# m1_3935_8137# sky130_fd_pr__res_xhigh_po_1p41_H3F4MM
Xsky130_fd_pr__nfet_g5v0d10v5_SB5CJ8_0 avss avss m1_10901_199# ena sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
C0 m1_179_3223# avss 0.217064f
C1 m1_179_5491# m1_179_6247# 0.011612f
C2 m1_3935_9649# m1_3935_10405# 0.011612f
C4 out_1010 out_1100 0.381021f
C5 m1_10911_14185# avss 0.217063f
C6 m1_179_7003# m1_179_6247# 0.011612f
C7 m1_7155_13051# m1_7155_12295# 0.011612f
C8 m1_179_2467# m1_179_1711# 0.011612f
C9 m1_179_3979# m1_179_4735# 0.011612f
C10 out_1011 out_1100 0.803817f
C11 m1_7155_1711# m1_7155_1333# 0.054565f
C12 m1_3399_8893# m1_3399_8137# 0.011612f
C13 m1_7155_2467# m1_7155_2845# 0.054566f
C14 m1_7155_9271# m1_7155_8515# 0.011612f
C15 m1_179_955# avss 0.216188f
C16 m1_179_8515# avss 0.217064f
C17 m1_3399_13429# m1_3935_13429# 0.044575f
C18 out_0100 out_0011 0.803817f
C19 out_0110 out_0111 0.280049f
C21 m1_3399_15697# m1_3399_16453# 0.011612f
C22 out_0100 m1_7155_8515# 0.083303f
C23 out_0110 out_0101 1.4187f
C24 m1_10901_8137# out_0110 0.013301f
C25 m1_3399_6625# m1_3935_6625# 0.044576f
C26 m1_7691_13807# m1_7691_13051# 0.011612f
C27 out_1111 m1_10911_2845# 0.071926f
C28 m1_10911_577# avss 0.214802f
C29 51 m1_7691_12295# 0.011612f
C30 avss m1_179_199# 0.092917f
C31 out_1000 m1_7691_7003# 0.020211f
C32 m1_3399_955# m1_3399_577# 0.054565f
C33 m1_179_11539# avss 0.217064f
C34 m1_179_6247# avss 0.217064f
C35 m1_3935_16453# m1_3935_15697# 0.011612f
C36 ena m1_10901_199# 0.333946f
C37 m1_10911_13429# m1_10911_14185# 0.011612f
C38 m1_179_14563# avss 0.217064f
C39 m1_3935_8137# m1_3399_8137# 0.044576f
C40 m1_10911_12673# avss 0.217063f
C41 m1_7155_7003# m1_7155_6247# 0.011612f
C42 m1_179_5491# m1_179_4735# 0.011612f
C43 m1_10911_12673# m1_10911_11917# 0.011612f
C44 out_1010 m1_7155_5491# 0.083303f
C45 m1_179_15319# avss 0.217064f
C46 m1_7691_15319# m1_7691_16075# 0.011612f
C47 m1_179_1711# avss 0.217064f
C48 out_0001 out_0000 0.280049f
C49 m1_3935_13429# m1_3935_14185# 0.011612f
C50 m1_179_13807# avss 0.217063f
C51 out_1001 out_0111 0.016886f
C52 m1_7155_7759# m1_7155_8515# 0.011612f
C53 m1_179_10027# avss 0.217064f
C54 m1_3935_9649# m1_3399_9649# 0.044576f
C55 m1_7155_2089# m1_7155_2467# 0.054565f
C56 m1_7691_9271# m1_7691_10027# 0.011612f
C57 m1_7155_11539# 51 0.044576f
C58 m1_7155_10027# m1_7691_10027# 0.044576f
C59 avdd m1_10911_16453# 0.077925f
C60 out_1101 avss 0.216735f
C61 m1_3399_6625# m1_3399_7381# 0.011612f
C62 m1_7155_13807# m1_7155_13051# 0.011612f
C63 m1_3399_8893# m1_3399_9649# 0.011612f
C64 m1_179_16831# m1_179_16075# 0.011612f
C65 m1_3935_5869# m1_3935_5113# 0.011612f
C66 m1_10911_12673# m1_10911_13429# 0.011612f
C67 m1_7155_6247# m1_7155_5491# 0.011612f
C68 out_1000 out_1010 0.381021f
C69 avss m1_179_4735# 0.217064f
C70 m1_3399_11161# m1_3399_10405# 0.011612f
C71 m1_179_955# m1_179_199# 0.011612f
C72 m1_179_13051# avss 0.217064f
C73 m1_10911_577# m1_10901_199# 0.071926f
C74 out_0111 avss 0.216736f
C75 m1_179_7003# m1_179_7759# 0.011612f
C76 m1_7691_16075# m1_7155_16831# 0.011612f
C77 avss out_0000 0.216735f
C79 m1_10901_8137# avss 0.217046f
C80 m1_10911_11917# out_0000 0.020211f
C81 m1_3399_15697# m1_3935_15697# 0.044576f
C82 m1_10911_1333# m1_10911_2089# 0.011612f
C83 m1_7155_16831# m1_7155_17209# 0.054565f
C84 m1_3399_15697# m1_3399_14941# 0.011612f
C85 m1_10911_2845# m1_10911_2089# 0.011612f
C86 m1_179_955# m1_179_1711# 0.011612f
C87 m1_3935_9649# m1_3935_8893# 0.011612f
C88 m1_3399_14185# m1_3399_13429# 0.011612f
C89 m1_7691_16075# m1_7155_16075# 0.044576f
C90 out_0100 out_0101 0.593278f
C91 m1_10901_8137# out_0100 0.671846f
C92 out_1111 avss 0.216735f
C93 m1_7691_9271# m1_7155_9271# 0.044576f
C94 out_1000 m1_7155_6247# 0.083303f
C95 m1_7155_9271# m1_7155_10027# 0.011612f
C96 m1_179_7759# avss 0.217063f
C97 m1_3399_5869# m1_3935_5869# 0.044576f
C98 m1_7691_9271# out_0100 0.020211f
C99 m1_7155_3979# m1_7155_4735# 0.011612f
C100 m1_3399_8893# m1_3935_8893# 0.044576f
C101 m1_3399_2845# m1_3399_3223# 0.054565f
C102 m1_7155_3979# out_1110 0.083303f
C103 out_1000 out_1001 1.4187f
C104 m1_179_15319# m1_179_14563# 0.011612f
C105 m1_10901_8137# out_0011 0.016875f
C106 m1_7691_15319# m1_7155_15319# 0.044576f
C107 m1_3399_3979# m1_3399_3601# 0.054565f
C108 out_1010 out_1011 1.4187f
C109 m1_7155_3601# out_1110 0.066858f
C110 m1_179_14563# m1_179_13807# 0.011612f
C111 m1_179_16075# avss 0.216189f
C112 m1_10911_15697# m1_10911_16453# 0.011612f
C113 m1_179_10783# avss 0.217063f
C114 m1_3935_11917# m1_3399_11917# 0.044576f
C115 m1_3935_7381# m1_3935_6625# 0.011612f
C116 out_0010 out_0001 0.280049f
C117 m1_7155_199# m1_7155_577# 0.054565f
C118 avss m1_10911_16453# 0.214804f
C119 m1_3935_10405# m1_3935_11161# 0.011612f
C120 m1_3399_14185# m1_3399_14941# 0.011612f
C121 m1_3399_3979# m1_3399_4357# 0.011612f
C122 m1_7155_7759# m1_7155_7003# 0.011612f
C123 m1_7691_13051# m1_7691_12295# 0.011612f
C124 m1_7155_7759# out_0101 0.083302f
C125 m1_3399_14185# m1_3935_14185# 0.044576f
C126 m1_179_12295# avss 0.217063f
C127 m1_3935_8137# m1_3935_8893# 0.011612f
C128 m1_3399_12673# m1_3399_11917# 0.011612f
C129 m1_3399_11161# m1_3399_11917# 0.011612f
C130 m1_3399_3601# m1_3399_3223# 0.054565f
C131 m1_7155_10783# m1_7691_10783# 0.044576f
C132 m1_7691_15319# m1_7691_14563# 0.011612f
C134 m1_3935_15697# m1_3935_14941# 0.011612f
C135 m1_179_8515# m1_179_7759# 0.011612f
C136 m1_3935_6625# m1_3935_5869# 0.011612f
C137 m1_3935_12673# m1_3935_11917# 0.011612f
C138 out_0010 avss 0.216735f
C139 out_1001 out_1010 0.803817f
C140 out_1001 out_1011 0.016886f
C141 m1_3399_14941# m1_3935_14941# 0.044576f
C142 m1_7155_16831# m1_7155_16075# 0.011612f
C143 out_1101 out_1100 1.4187f
C144 m1_179_13051# m1_179_13807# 0.011612f
C145 m1_3399_4357# m1_3399_5113# 0.011612f
C146 m1_3935_14941# m1_3935_14185# 0.011612f
C147 m1_10911_1333# avss 0.217022f
C148 m1_3399_7381# m1_3935_7381# 0.044576f
C149 m1_7155_16075# m1_7155_15319# 0.011612f
C150 m1_3935_12673# m1_3399_12673# 0.044576f
C151 m1_7691_13807# m1_7155_13807# 0.044576f
C152 avss m1_10911_2089# 0.217063f
C153 m1_10911_2845# avss 0.217063f
C154 m1_3935_5113# m1_3399_5113# 0.044576f
C155 m1_3399_4357# m1_3935_4357# 0.044576f
C157 m1_179_3979# avss 0.217063f
C158 m1_3399_1333# m1_3399_955# 0.054565f
C159 out_0110 avss 0.216735f
C160 out_1011 avss 0.216735f
C161 m1_179_9271# avss 0.217063f
C162 m1_179_11539# m1_179_10783# 0.011612f
C163 out_0010 out_0011 0.280049f
C164 m1_3399_1711# m1_3399_2089# 0.054565f
C165 m1_3935_4357# m1_3935_5113# 0.011612f
C166 m1_179_16831# avss 0.092918f
C167 m1_3935_12673# m1_3935_13429# 0.011612f
C168 m1_7155_3601# m1_7155_3223# 0.054565f
C169 out_1101 out_1111 0.016886f
C170 m1_10901_8137# out_0101 0.058289f
C171 m1_7691_13051# m1_7155_13051# 0.044576f
C172 m1_179_11539# m1_179_12295# 0.011612f
C173 m1_179_15319# m1_179_16075# 0.011612f
C174 m1_3399_2089# m1_3399_2467# 0.054565f
C175 m1_179_2467# avss 0.217063f
C176 m1_179_10783# m1_179_10027# 0.011612f
C177 m1_3399_5869# m1_3399_5113# 0.011612f
C178 m1_3399_10405# m1_3935_10405# 0.044576f
C179 m1_7691_13807# m1_7691_14563# 0.011612f
C180 m1_3935_8137# m1_3935_7381# 0.011612f
C181 m1_179_3979# m1_179_3223# 0.011612f
C182 out_0001 avss 0.216735f
C183 m1_179_5491# avss 0.217063f
C184 m1_7155_10783# m1_7155_11539# 0.011612f
C185 m1_7155_12295# m1_7691_12295# 0.044576f
C186 m1_7155_10783# m1_7155_10027# 0.011612f
C187 m1_7155_3601# m1_7155_3979# 0.011612f
C188 out_1101 out_1110 0.803817f
C189 out_1001 avss 0.216735f
C190 m1_179_7003# avss 0.217064f
C191 m1_7155_955# m1_7155_1333# 0.054565f
C192 m1_10911_577# m1_10911_1333# 0.011612f
C193 m1_3399_2845# m1_3399_2467# 0.054565f
C194 m1_7155_4735# out_1100 0.083303f
C195 m1_7155_3223# m1_7155_2845# 0.054565f
C196 m1_7155_955# m1_7155_577# 0.054565f
C197 m1_10911_14941# m1_10911_15697# 0.011612f
C198 out_1110 out_1100 0.381021f
C199 m1_179_8515# m1_179_9271# 0.011612f
C200 m1_7155_13807# m1_7155_14563# 0.011612f
C201 m1_10911_14941# avss 0.217063f
C202 m1_179_2467# m1_179_3223# 0.011612f
C203 m1_7155_1711# m1_7155_2089# 0.054565f
C204 m1_10911_15697# avss 0.217022f
C205 m1_179_12295# m1_179_13051# 0.011612f
C206 m1_3399_3979# m1_3935_4357# 0.011612f
C207 m1_3399_16453# m1_3935_16453# 0.044576f
C208 m1_7155_11539# m1_7155_12295# 0.011612f
C209 out_1000 out_0111 0.803817f
C210 m1_3399_6625# m1_3399_5869# 0.011612f
C211 m1_7155_14563# m1_7155_15319# 0.011612f
C212 m1_7155_7003# m1_7691_7003# 0.044576f
C213 m1_10911_11917# avss 0.217064f
C214 out_1000 out_0101 0.129936f
C215 out_0101 m1_7691_7003# 0.071926f
C216 m1_3935_11917# m1_3935_11161# 0.011612f
C217 m1_7691_10783# m1_7691_10027# 0.011612f
C218 out_1111 out_1110 1.4187f
C219 m1_3399_10405# m1_3399_9649# 0.011612f
C220 m1_7691_10783# 51 0.011612f
C222 m1_7155_5491# m1_7155_4735# 0.011612f
C223 m1_3399_16453# m1_3399_17209# 0.011612f
C224 m1_3399_11161# m1_3935_11161# 0.044576f
C225 m1_179_9271# m1_179_10027# 0.011612f
C226 m1_3399_7381# m1_3399_8137# 0.011612f
C228 m1_3399_13429# m1_3399_12673# 0.011612f
C229 m1_10911_14941# m1_10911_14185# 0.011612f
C230 m1_3399_17209# m1_3935_16453# 0.011612f
C231 m1_3399_1711# m1_3399_1333# 0.054565f
C232 m1_3399_199# m1_3399_577# 0.054565f
C233 out_1101 out_1011 0.016886f
C234 m1_10911_13429# avss 0.217063f
C235 m1_7691_14563# m1_7155_14563# 0.044576f
C236 out_0011 avss 0.216735f
C237 ena 0 3.253165f
C238 avdd 0 8.495175f
C239 m1_10911_16453# 0 0.789952f
C240 m1_7691_16075# 0 0.600369f
C241 m1_10911_15697# 0 0.789096f
C242 m1_7691_15319# 0 0.599493f
C243 m1_10911_14941# 0 0.789055f
C244 m1_7691_14563# 0 0.599493f
C245 m1_10911_14185# 0 0.789055f
C246 m1_7691_13807# 0 0.599493f
C247 m1_10911_13429# 0 0.789055f
C248 m1_7691_13051# 0 0.599493f
C249 m1_10911_12673# 0 0.789055f
C250 m1_7691_12295# 0 0.599493f
C251 m1_10911_11917# 0 0.789055f
C252 51 0 0.599493f
C253 out_0000 0 3.014127f
C254 out_0001 0 2.851987f
C255 m1_7691_10783# 0 0.599493f
C256 m1_7691_10027# 0 0.599493f
C257 out_0010 0 2.851987f
C258 out_0011 0 2.656507f
C259 m1_7691_9271# 0 0.599493f
C260 out_0100 0 2.947894f
C261 m1_10901_8137# 0 0.800173f
C262 out_0110 0 2.696149f
C263 out_0101 0 2.833084f
C264 out_0111 0 2.656507f
C265 m1_7691_7003# 0 0.599493f
C266 out_1001 0 2.500679f
C267 out_1000 0 2.668634f
C268 out_1011 0 2.500679f
C269 out_1010 0 2.564904f
C270 out_1101 0 2.500679f
C271 out_1100 0 2.564904f
C272 out_1111 0 2.860089f
C273 out_1110 0 2.790774f
C274 m1_10911_2845# 0 0.789055f
C275 m1_10911_2089# 0 0.789055f
C276 m1_10911_1333# 0 0.789096f
C277 m1_10911_577# 0 0.791315f
C278 m1_10901_199# 0 3.463708f
C279 m1_7155_17209# 0 0.883249f
C280 m1_7155_16831# 0 0.604193f
C281 m1_3935_16453# 0 0.601754f
C282 m1_7155_16075# 0 0.600369f
C283 m1_3935_15697# 0 0.599535f
C284 m1_7155_15319# 0 0.599493f
C285 m1_3935_14941# 0 0.599493f
C286 m1_7155_14563# 0 0.599493f
C287 m1_3935_14185# 0 0.599493f
C288 m1_7155_13807# 0 0.599493f
C289 m1_3935_13429# 0 0.599493f
C290 m1_7155_13051# 0 0.599493f
C291 m1_3935_12673# 0 0.599493f
C292 m1_7155_12295# 0 0.599493f
C293 m1_3935_11917# 0 0.599493f
C294 m1_7155_11539# 0 0.599493f
C295 m1_3935_11161# 0 0.599493f
C296 m1_7155_10783# 0 0.599493f
C297 m1_3935_10405# 0 0.599493f
C298 m1_7155_10027# 0 0.599493f
C299 m1_3935_9649# 0 0.599493f
C300 m1_7155_9271# 0 0.599493f
C301 m1_3935_8893# 0 0.599493f
C302 m1_7155_8515# 0 0.598612f
C303 m1_3935_8137# 0 0.599493f
C304 m1_7155_7759# 0 0.598612f
C305 m1_3935_7381# 0 0.599493f
C306 m1_7155_7003# 0 0.599493f
C307 m1_3935_6625# 0 0.599493f
C308 m1_7155_6247# 0 0.598612f
C309 m1_3935_5869# 0 0.599493f
C310 m1_7155_5491# 0 0.598612f
C311 m1_3935_5113# 0 0.599493f
C312 m1_7155_4735# 0 0.598612f
C313 m1_3935_4357# 0 0.599493f
C314 m1_7155_3979# 0 0.598612f
C315 m1_7155_3601# 0 0.599576f
C316 m1_7155_3223# 0 0.583453f
C317 m1_7155_2845# 0 0.583453f
C318 m1_7155_2467# 0 0.583453f
C319 m1_7155_2089# 0 0.583453f
C320 m1_7155_1711# 0 0.583453f
C321 m1_7155_1333# 0 0.583545f
C322 m1_7155_955# 0 0.584937f
C323 m1_7155_577# 0 0.586355f
C324 m1_7155_199# 0 0.883249f
C325 m1_3399_17209# 0 0.901087f
C326 m1_179_16831# 0 0.924812f
C327 m1_3399_16453# 0 0.601754f
C328 m1_179_16075# 0 0.78993f
C329 m1_3399_15697# 0 0.599535f
C330 m1_179_15319# 0 0.789055f
C331 m1_3399_14941# 0 0.599493f
C332 m1_179_14563# 0 0.789055f
C333 m1_3399_14185# 0 0.599493f
C334 m1_179_13807# 0 0.789055f
C335 m1_3399_13429# 0 0.599493f
C336 m1_179_13051# 0 0.789055f
C337 m1_3399_12673# 0 0.599493f
C338 m1_179_12295# 0 0.789055f
C339 m1_3399_11917# 0 0.599493f
C340 m1_179_11539# 0 0.789055f
C341 m1_3399_11161# 0 0.599493f
C342 m1_179_10783# 0 0.789055f
C343 m1_3399_10405# 0 0.599493f
C344 m1_179_10027# 0 0.789055f
C345 m1_3399_9649# 0 0.599493f
C346 m1_179_9271# 0 0.789055f
C347 m1_3399_8893# 0 0.599493f
C348 m1_179_8515# 0 0.789055f
C349 m1_3399_8137# 0 0.599493f
C350 m1_179_7759# 0 0.789055f
C351 m1_3399_7381# 0 0.599493f
C352 m1_179_7003# 0 0.789055f
C353 m1_3399_6625# 0 0.599493f
C354 m1_179_6247# 0 0.789055f
C355 m1_3399_5869# 0 0.599493f
C356 m1_179_5491# 0 0.789055f
C357 m1_3399_5113# 0 0.599493f
C358 m1_179_4735# 0 0.789055f
C359 m1_3399_4357# 0 0.599493f
C360 m1_3399_3979# 0 0.601291f
C361 m1_179_3979# 0 0.789055f
C362 m1_3399_3601# 0 0.583453f
C363 m1_3399_3223# 0 0.583453f
C364 m1_179_3223# 0 0.789055f
C365 m1_3399_2845# 0 0.583453f
C366 m1_3399_2467# 0 0.583453f
C367 m1_179_2467# 0 0.789055f
C368 m1_3399_2089# 0 0.583453f
C369 m1_3399_1711# 0 0.583453f
C370 m1_179_1711# 0 0.789055f
C371 m1_3399_1333# 0 0.583545f
C372 m1_3399_955# 0 0.584937f
C373 m1_179_955# 0 0.78993f
C374 m1_3399_577# 0 0.586355f
C375 m1_3399_199# 0 0.883249f
C376 m1_179_199# 0 0.924812f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100# 0
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 w_n558_n397# a_300_n100# 0.081002f
C1 a_n300_n197# w_n558_n397# 1.02259f
C2 a_n300_n197# a_300_n100# 0.042408f
C3 w_n558_n397# a_n358_n100# 0.081002f
C4 a_n358_n100# a_300_n100# 0.021684f
C5 a_n300_n197# a_n358_n100# 0.042408f
C6 a_300_n100# 0 0.067884f
C7 a_n358_n100# 0 0.067884f
C8 a_n300_n197# 0 0.770863f
C9 w_n558_n397# 0 3.43953f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CY564Z a_300_n100# a_n492_n322# a_n358_n100#
+ a_n300_n188#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n492_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 a_n358_n100# a_n300_n188# 0.042408f
C1 a_n300_n188# a_300_n100# 0.042408f
C2 a_n358_n100# a_300_n100# 0.021684f
C3 a_300_n100# a_n492_n322# 0.148584f
C4 a_n358_n100# a_n492_n322# 0.148584f
C5 a_n300_n188# a_n492_n322# 1.74754f
.ends

.subckt trans_gate_m in ena_b ena out avdd vss
Xsky130_fd_pr__pfet_g5v0d10v5_6H9SQ3_1 ena_b out avdd in vss sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3
Xsky130_fd_pr__nfet_g5v0d10v5_CY564Z_0 out vss in ena sky130_fd_pr__nfet_g5v0d10v5_CY564Z
C0 avdd out 0.092004f
C1 ena_b avdd 0.220595f
C2 ena_b out 0.095084f
C3 avdd in 0.379728f
C4 avdd ena 0.070299f
C5 in out 0.018089f
C6 ena out 0.092409f
C7 ena_b in 0.095084f
C8 ena_b ena 0.066395f
C9 ena in 0.092409f
C10 ena vss 1.902743f
C11 out vss 0.619585f
C12 in vss 0.331515f
C13 ena_b vss 0.779553f
C14 avdd vss 4.054391f
.ends

.subckt multiplexer in_0000 in_0001 in_0011 in_0100 in_0101 in_0110 vtrip_3 vtrip_3_b
+ vtrip_2 out vtrip_1_b in_1000 in_1001 in_1010 in_1100 in_1101 in_1110 in_1111 trans_gate_m_37/in
+ trans_gate_m_32/in vtrip_0_b trans_gate_m_7/out in_1011 trans_gate_m_27/in trans_gate_m_3/out
+ trans_gate_m_33/in trans_gate_m_34/in trans_gate_m_28/in in_0111 in_0010 trans_gate_m_5/out
+ trans_gate_m_20/in trans_gate_m_31/in trans_gate_m_23/in trans_gate_m_9/out vtrip_2_b
+ trans_gate_m_29/in vss vtrip_1 vtrip_0 avdd
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_2 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_3 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_4 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_5 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_6 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_7 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_8 vss vtrip_2_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_9 vss vtrip_2 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_20 trans_gate_m_20/in vtrip_2 vtrip_2_b trans_gate_m_33/in avdd vss
+ trans_gate_m
Xtrans_gate_m_31 trans_gate_m_31/in vtrip_1 vtrip_1_b trans_gate_m_20/in avdd vss
+ trans_gate_m
Xtrans_gate_m_0 in_0010 vtrip_0 vtrip_0_b trans_gate_m_29/in avdd vss trans_gate_m
Xtrans_gate_m_1 in_0011 vtrip_0_b vtrip_0 trans_gate_m_29/in avdd vss trans_gate_m
Xtrans_gate_m_10 in_1000 vtrip_0 vtrip_0_b trans_gate_m_23/in avdd vss trans_gate_m
Xtrans_gate_m_21 trans_gate_m_5/out vtrip_1_b vtrip_1 trans_gate_m_32/in avdd vss
+ trans_gate_m
Xtrans_gate_m_32 trans_gate_m_32/in vtrip_2 vtrip_2_b trans_gate_m_34/in avdd vss
+ trans_gate_m
Xtrans_gate_m_2 in_0110 vtrip_0 vtrip_0_b trans_gate_m_3/out avdd vss trans_gate_m
Xtrans_gate_m_11 in_1001 vtrip_0_b vtrip_0 trans_gate_m_23/in avdd vss trans_gate_m
Xtrans_gate_m_33 trans_gate_m_33/in vtrip_3 vtrip_3_b out avdd vss trans_gate_m
Xtrans_gate_m_3 in_0111 vtrip_0_b vtrip_0 trans_gate_m_3/out avdd vss trans_gate_m
Xtrans_gate_m_12 in_0101 vtrip_0_b vtrip_0 trans_gate_m_27/in avdd vss trans_gate_m
Xtrans_gate_m_23 trans_gate_m_23/in vtrip_1 vtrip_1_b trans_gate_m_32/in avdd vss
+ trans_gate_m
Xtrans_gate_m_34 trans_gate_m_34/in vtrip_3_b vtrip_3 out avdd vss trans_gate_m
Xtrans_gate_m_4 in_1011 vtrip_0_b vtrip_0 trans_gate_m_5/out avdd vss trans_gate_m
Xtrans_gate_m_13 in_0100 vtrip_0 vtrip_0_b trans_gate_m_27/in avdd vss trans_gate_m
Xtrans_gate_m_5 in_1010 vtrip_0 vtrip_0_b trans_gate_m_5/out avdd vss trans_gate_m
Xtrans_gate_m_14 in_0001 vtrip_0_b vtrip_0 trans_gate_m_31/in avdd vss trans_gate_m
Xtrans_gate_m_25 trans_gate_m_3/out vtrip_1_b vtrip_1 trans_gate_m_28/in avdd vss
+ trans_gate_m
Xtrans_gate_m_6 in_1110 vtrip_0 vtrip_0_b trans_gate_m_7/out avdd vss trans_gate_m
Xtrans_gate_m_15 in_0000 vtrip_0 vtrip_0_b trans_gate_m_31/in avdd vss trans_gate_m
Xtrans_gate_m_27 trans_gate_m_27/in vtrip_1 vtrip_1_b trans_gate_m_28/in avdd vss
+ trans_gate_m
Xtrans_gate_m_37 trans_gate_m_37/in vtrip_2_b vtrip_2 trans_gate_m_34/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_10 vss vtrip_3_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_7 in_1111 vtrip_0_b vtrip_0 trans_gate_m_7/out avdd vss trans_gate_m
Xtrans_gate_m_28 trans_gate_m_28/in vtrip_2_b vtrip_2 trans_gate_m_33/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_11 vss vtrip_3 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_8 in_1101 vtrip_0_b vtrip_0 trans_gate_m_9/out avdd vss trans_gate_m
Xtrans_gate_m_18 trans_gate_m_9/out vtrip_1 vtrip_1_b trans_gate_m_37/in avdd vss
+ trans_gate_m
Xtrans_gate_m_29 trans_gate_m_29/in vtrip_1_b vtrip_1 trans_gate_m_20/in avdd vss
+ trans_gate_m
Xtrans_gate_m_9 in_1100 vtrip_0 vtrip_0_b trans_gate_m_9/out avdd vss trans_gate_m
Xtrans_gate_m_19 trans_gate_m_7/out vtrip_1_b vtrip_1 trans_gate_m_37/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_1 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
C0 in_1011 vtrip_0_b 0.303747f
C1 trans_gate_m_7/out vtrip_0_b 0.015828f
C2 in_1111 vtrip_0 0.085069f
C3 in_0011 trans_gate_m_31/in 0.183189f
C4 in_1111 trans_gate_m_9/out 0.183189f
C5 in_1110 vtrip_0 0.10236f
C6 trans_gate_m_29/in trans_gate_m_27/in 0.010259f
C7 in_1110 trans_gate_m_9/out 0.204661f
C8 trans_gate_m_3/out trans_gate_m_23/in 0.010259f
C9 trans_gate_m_7/out vtrip_1 0.828205f
C10 trans_gate_m_28/in vtrip_2 0.883815f
C11 in_0011 vtrip_0 0.10287f
C12 trans_gate_m_5/out trans_gate_m_23/in 0.362471f
C13 trans_gate_m_28/in vtrip_2_b 0.466992f
C14 trans_gate_m_27/in in_0111 0.183189f
C15 trans_gate_m_27/in in_0110 0.204661f
C16 in_0111 in_1010 0.144733f
C17 trans_gate_m_5/out trans_gate_m_9/out 0.010259f
C18 vtrip_2 trans_gate_m_20/in 0.612399f
C19 vtrip_2_b trans_gate_m_20/in 0.318836f
C20 avdd trans_gate_m_23/in 0.345067f
C21 trans_gate_m_31/in avdd 0.341363f
C22 in_1000 in_1010 0.044575f
C23 trans_gate_m_37/in vtrip_2 0.551211f
C24 in_0010 in_0000 0.044575f
C25 in_0110 in_0111 0.098921f
C26 trans_gate_m_37/in vtrip_2_b 0.309159f
C27 in_1111 in_1101 0.044575f
C28 avdd vtrip_0 8.880435f
C29 trans_gate_m_28/in avdd 0.235617f
C30 in_1111 vtrip_0_b 0.321101f
C31 avdd trans_gate_m_9/out 0.341586f
C32 vtrip_0_b in_1110 0.303873f
C33 in_1100 in_1001 0.026216f
C34 in_0011 vtrip_0_b 0.303747f
C35 trans_gate_m_7/out vtrip_1_b 0.424647f
C36 trans_gate_m_32/in vtrip_2 0.901041f
C37 trans_gate_m_20/in avdd 0.229713f
C38 trans_gate_m_32/in vtrip_2_b 0.443648f
C39 trans_gate_m_3/out vtrip_0_b 0.015722f
C40 vtrip_1 vtrip_2 0.01408f
C41 trans_gate_m_5/out vtrip_0_b 0.015722f
C42 trans_gate_m_37/in avdd 0.212793f
C43 vtrip_1 vtrip_2_b 0.165901f
C44 avdd in_1001 0.186342f
C45 in_1100 in_1101 0.026216f
C46 trans_gate_m_3/out vtrip_1 0.827916f
C47 vtrip_3 trans_gate_m_33/in 0.531277f
C48 in_1011 in_1010 0.098921f
C49 vtrip_1 trans_gate_m_5/out 0.827916f
C50 vtrip_3 vtrip_2_b 0.015168f
C51 in_0101 in_0100 0.026216f
C52 in_1101 avdd 0.175548f
C53 avdd vtrip_0_b 2.747238f
C54 trans_gate_m_32/in avdd 0.220392f
C55 trans_gate_m_23/in vtrip_0 1.164039f
C56 trans_gate_m_31/in vtrip_0 1.154617f
C57 vtrip_3 vtrip_3_b 0.90924f
C58 trans_gate_m_23/in trans_gate_m_9/out 0.011864f
C59 vtrip_1 avdd 8.547259f
C60 in_0100 avdd 0.186342f
C61 trans_gate_m_9/out vtrip_0 1.154381f
C62 vtrip_3 avdd 2.240629f
C63 in_0001 in_0100 0.026216f
C64 trans_gate_m_31/in trans_gate_m_20/in 0.011995f
C65 vtrip_2 vtrip_1_b 0.017624f
C66 vtrip_2_b vtrip_1_b 0.603929f
C67 trans_gate_m_3/out vtrip_1_b 0.332586f
C68 trans_gate_m_28/in trans_gate_m_20/in 0.033198f
C69 trans_gate_m_5/out vtrip_1_b 0.332586f
C70 trans_gate_m_37/in trans_gate_m_9/out 0.013606f
C71 in_0011 trans_gate_m_29/in 0.013238f
C72 trans_gate_m_23/in vtrip_0_b 1.297016f
C73 trans_gate_m_31/in vtrip_0_b 1.401507f
C74 trans_gate_m_3/out trans_gate_m_27/in 0.362471f
C75 trans_gate_m_3/out trans_gate_m_29/in 0.033198f
C76 trans_gate_m_32/in trans_gate_m_23/in 0.013606f
C77 avdd in_0000 0.185437f
C78 avdd vtrip_1_b 2.36787f
C79 vtrip_1 trans_gate_m_23/in 0.043456f
C80 vtrip_0_b vtrip_0 3.714523f
C81 vtrip_1 trans_gate_m_31/in 0.040929f
C82 in_0011 in_0110 0.144733f
C83 in_0001 in_0000 0.026216f
C84 vtrip_0_b trans_gate_m_9/out 1.405763f
C85 trans_gate_m_28/in trans_gate_m_32/in 0.031058f
C86 trans_gate_m_3/out in_0111 0.013238f
C87 vtrip_1 vtrip_0 0.060603f
C88 vtrip_1 trans_gate_m_9/out 0.043808f
C89 in_0101 in_0111 0.044575f
C90 trans_gate_m_27/in avdd 0.345558f
C91 trans_gate_m_33/in trans_gate_m_34/in 0.031154f
C92 in_1010 avdd 0.181177f
C93 trans_gate_m_29/in avdd 0.235334f
C94 vtrip_2_b trans_gate_m_34/in 0.029424f
C95 in_1000 in_0101 0.026216f
C96 trans_gate_m_32/in trans_gate_m_37/in 0.033198f
C97 in_0111 avdd 0.189004f
C98 in_0110 avdd 0.181177f
C99 in_0011 in_0010 0.098921f
C100 vtrip_3_b trans_gate_m_34/in 0.319358f
C101 in_1000 avdd 0.186342f
C102 trans_gate_m_7/out in_1111 0.013238f
C103 trans_gate_m_23/in vtrip_1_b 0.738587f
C104 trans_gate_m_31/in vtrip_1_b 0.786715f
C105 in_1011 in_1110 0.144733f
C106 avdd trans_gate_m_34/in 0.197834f
C107 vtrip_0 vtrip_1_b 0.210797f
C108 trans_gate_m_28/in vtrip_1_b 0.021556f
C109 trans_gate_m_9/out vtrip_1_b 0.74635f
C110 trans_gate_m_5/out in_1011 0.013238f
C111 trans_gate_m_7/out trans_gate_m_5/out 0.033198f
C112 trans_gate_m_27/in trans_gate_m_23/in 0.011864f
C113 trans_gate_m_27/in trans_gate_m_31/in 0.011864f
C114 in_1010 trans_gate_m_23/in 0.204661f
C115 trans_gate_m_29/in trans_gate_m_31/in 0.36247f
C116 avdd in_0010 0.173735f
C117 trans_gate_m_20/in vtrip_1_b 0.021662f
C118 trans_gate_m_27/in vtrip_0 1.155297f
C119 trans_gate_m_28/in trans_gate_m_27/in 0.011995f
C120 in_1010 vtrip_0 0.10236f
C121 trans_gate_m_37/in vtrip_1_b 0.021592f
C122 in_1011 avdd 0.189004f
C123 trans_gate_m_7/out avdd 0.22238f
C124 in_0111 vtrip_0 0.10287f
C125 in_0110 vtrip_0 0.10001f
C126 in_1111 in_1110 0.098921f
C127 vtrip_0_b vtrip_1_b 0.557411f
C128 trans_gate_m_32/in vtrip_1_b 0.021486f
C129 vtrip_2 vtrip_2_b 2.141323f
C130 vtrip_1 vtrip_1_b 3.174343f
C131 trans_gate_m_33/in vtrip_2_b 0.029429f
C132 out vtrip_3_b 0.023178f
C133 trans_gate_m_31/in in_0010 0.204661f
C134 trans_gate_m_27/in vtrip_0_b 1.297017f
C135 trans_gate_m_29/in vtrip_0_b 0.015828f
C136 in_1100 in_1110 0.044575f
C137 in_1010 vtrip_0_b 0.303873f
C138 out avdd 0.050125f
C139 vtrip_2 vtrip_3_b 0.061436f
C140 trans_gate_m_33/in vtrip_3_b 0.338688f
C141 in_1000 in_1001 0.026216f
C142 trans_gate_m_3/out trans_gate_m_5/out 0.033198f
C143 in_0010 vtrip_0 0.086196f
C144 vtrip_1 trans_gate_m_27/in 0.041106f
C145 in_1111 avdd 0.143003f
C146 vtrip_3_b vtrip_2_b 0.210613f
C147 vtrip_1 trans_gate_m_29/in 0.827921f
C148 in_1011 trans_gate_m_23/in 0.183189f
C149 avdd in_1110 0.181177f
C150 in_0111 vtrip_0_b 0.303747f
C151 in_0110 vtrip_0_b 0.303873f
C152 vtrip_2 avdd 6.213146f
C153 trans_gate_m_33/in avdd 0.233559f
C154 in_0011 avdd 0.189004f
C155 in_1011 vtrip_0 0.10287f
C156 vtrip_2_b avdd 1.632203f
C157 trans_gate_m_7/out trans_gate_m_9/out 0.362471f
C158 trans_gate_m_3/out avdd 0.235333f
C159 in_0011 in_0001 0.044575f
C160 in_0110 in_0100 0.044575f
C161 trans_gate_m_5/out avdd 0.235334f
C162 in_0101 avdd 0.186342f
C163 in_1100 avdd 0.186342f
C164 vtrip_3_b avdd 0.58496f
C165 in_1011 in_1001 0.044575f
C166 vtrip_0_b in_0010 0.320617f
C167 vtrip_3 trans_gate_m_34/in 0.594121f
C168 trans_gate_m_27/in vtrip_1_b 0.738587f
C169 trans_gate_m_29/in vtrip_1_b 0.383684f
C170 in_0001 avdd 0.186342f
C171 vtrip_1 vss 12.708198f
C172 in_1100 vss 0.331279f
C173 trans_gate_m_20/in vss 2.707844f
C174 vtrip_1_b vss 10.844804f
C175 trans_gate_m_37/in vss 2.744655f
C176 vtrip_0 vss 22.511623f
C177 trans_gate_m_9/out vss 3.423639f
C178 in_1101 vss 0.382099f
C179 vtrip_0_b vss 20.25898f
C180 trans_gate_m_33/in vss 4.255809f
C181 in_1111 vss 0.688102f
C182 vtrip_2 vss 7.108443f
C183 trans_gate_m_34/in vss 4.259955f
C184 vtrip_2_b vss 7.432176f
C185 avdd vss 0.113819p
C186 in_0000 vss 0.371548f
C187 trans_gate_m_7/out vss 2.612008f
C188 in_1110 vss 0.424785f
C189 trans_gate_m_28/in vss 2.5033f
C190 trans_gate_m_31/in vss 3.449917f
C191 in_0001 vss 0.331279f
C192 in_1010 vss 0.424785f
C193 in_0100 vss 0.331279f
C194 trans_gate_m_5/out vss 2.51077f
C195 in_1011 vss 0.425005f
C196 vtrip_3 vss 3.874589f
C197 out vss 2.697432f
C198 vtrip_3_b vss 3.233042f
C199 trans_gate_m_27/in vss 3.409393f
C200 in_0101 vss 0.331279f
C201 trans_gate_m_3/out vss 2.510769f
C202 in_0111 vss 0.425005f
C203 trans_gate_m_23/in vss 3.407793f
C204 in_1001 vss 0.331279f
C205 in_0110 vss 0.424785f
C206 trans_gate_m_32/in vss 2.509769f
C207 in_1000 vss 0.331279f
C208 trans_gate_m_29/in vss 2.592289f
C209 in_0011 vss 0.425005f
C210 in_0010 vss 0.647162f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YHAZV5 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100# 0
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 w_n558_n397# a_n300_n197# 1.02259f
C1 w_n558_n397# a_300_n100# 0.081002f
C2 a_300_n100# a_n300_n197# 0.042408f
C3 w_n558_n397# a_n358_n100# 0.081002f
C4 a_n300_n197# a_n358_n100# 0.042408f
C5 a_300_n100# a_n358_n100# 0.021684f
C6 a_300_n100# 0 0.067884f
C7 a_n358_n100# 0 0.067884f
C8 a_n300_n197# 0 0.770863f
C9 w_n558_n397# 0 3.43953f
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_37RBXE a_n147_n172# a_n45_n70#
X0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
C0 a_n45_n70# a_n147_n172# 0.219937f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EEVBR7 a_n300_n288# a_300_n200# a_n492_n422#
+ a_n358_n200#
X0 a_300_n200# a_n300_n288# a_n358_n200# a_n492_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
C0 a_n300_n288# a_n358_n200# 0.077833f
C1 a_n300_n288# a_300_n200# 0.077833f
C2 a_n358_n200# a_300_n200# 0.043012f
C3 a_300_n200# a_n492_n422# 0.265261f
C4 a_n358_n200# a_n492_n422# 0.265261f
C5 a_n300_n288# a_n492_n422# 1.78694f
.ends

.subckt sky130_fd_pr__nfet_01v8_MG6U6H a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 a_n300_n188# a_n358_n100# 0.042408f
C1 a_n300_n188# a_300_n100# 0.042408f
C2 a_n358_n100# a_300_n100# 0.021684f
C3 a_300_n100# a_n460_n274# 0.157496f
C4 a_n358_n100# a_n460_n274# 0.157496f
C5 a_n300_n188# a_n460_n274# 1.84766f
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9Q3 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 w_n496_n319# a_n300_n197# 1.05203f
C1 w_n496_n319# a_300_n100# 0.085201f
C2 a_300_n100# a_n300_n197# 0.042408f
C3 w_n496_n319# a_n358_n100# 0.085201f
C4 a_n300_n197# a_n358_n100# 0.042408f
C5 a_300_n100# a_n358_n100# 0.021684f
C6 a_300_n100# 0 0.071857f
C7 a_n358_n100# 0 0.071857f
C8 a_n300_n197# 0 0.838987f
C9 w_n496_n319# 0 2.60523f
.ends

.subckt level_shifter in out out_b dvss in_b avss M2 avdd
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0 out_b out avdd avdd avss sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1 out out_b avdd avdd avss sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__diode_pw2nd_05v5_37RBXE_0 dvss in sky130_fd_pr__diode_pw2nd_05v5_37RBXE
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0 in_b out avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1 in out_b avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_01v8_MG6U6H_0 dvss in_b in dvss sky130_fd_pr__nfet_01v8_MG6U6H
Xsky130_fd_pr__pfet_01v8_J2L9Q3_0 in in_b M2 M2 sky130_fd_pr__pfet_01v8_J2L9Q3
C0 avdd out_b 0.344028f
C1 out out_b 1.515421f
C2 avdd out 0.595998f
C3 in in_b 2.070184f
C4 in M2 0.777228f
C5 in dvss 1.323499f
C6 in_b M2 0.258043f
C7 in_b dvss 0.401345f
C8 dvss M2 5.414917f
C9 in out_b 0.080172f
C10 avdd in 0.023962f
C11 in out 0.035795f
C12 in_b out_b 0.073298f
C13 avdd in_b 0.018185f
C14 in_b out 0.077183f
C15 M2 sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 7.777787f
C16 dvss sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 0.08954f
C17 in sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 5.468968f
C18 in_b sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 3.504763f
C19 out_b sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 1.443518f
C20 out sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 1.328238f
C21 avdd sky130_fd_pr__pfet_01v8_J2L9Q3_0/0 7.069616f
.ends

.subckt sky130_fd_pr__pfet_01v8_XTWSDC a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
+ 0
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
C0 w_n1796_n319# a_n1658_n100# 0.085193f
C1 w_n1796_n319# a_n1600_n197# 5.05964f
C2 a_1600_n100# w_n1796_n319# 0.085193f
C3 a_n1658_n100# a_n1600_n197# 0.049339f
C4 a_1600_n100# a_n1600_n197# 0.049339f
C5 a_1600_n100# 0 0.091337f
C6 a_n1658_n100# 0 0.091337f
C7 a_n1600_n197# 0 4.27103f
C8 w_n1796_n319# 0 8.81803f
.ends

.subckt sky130_fd_pr__nfet_01v8_7ZF23Z a_2000_n100# a_n2058_n100# a_n2000_n188# a_n2160_n274#
X0 a_2000_n100# a_n2000_n188# a_n2058_n100# a_n2160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
C0 a_n2000_n188# a_2000_n100# 0.049339f
C1 a_n2000_n188# a_n2058_n100# 0.049339f
C2 a_2000_n100# a_n2160_n274# 0.176968f
C3 a_n2058_n100# a_n2160_n274# 0.176968f
C4 a_n2000_n188# a_n2160_n274# 11.3874f
.ends

.subckt sky130_fd_pr__nfet_01v8_V433WY a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 a_n300_n188# a_300_n100# 0.042408f
C1 a_n300_n188# a_n358_n100# 0.042408f
C2 a_300_n100# a_n358_n100# 0.021684f
C3 a_300_n100# a_n460_n274# 0.157496f
C4 a_n358_n100# a_n460_n274# 0.157496f
C5 a_n300_n188# a_n460_n274# 1.84766f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69BJMM a_n500_n188# a_500_n100# a_n692_n322#
+ a_n558_n100#
X0 a_500_n100# a_n500_n188# a_n558_n100# a_n692_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
C0 a_n500_n188# a_500_n100# 0.046765f
C1 a_n500_n188# a_n558_n100# 0.046765f
C2 a_500_n100# a_n558_n100# 0.013433f
C3 a_500_n100# a_n692_n322# 0.15299f
C4 a_n558_n100# a_n692_n322# 0.15299f
C5 a_n500_n188# a_n692_n322# 2.80683f
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E7V9VM w_n758_n897# a_n558_n600# a_n500_n697#
+ a_500_n600# 0
X0 a_500_n600# a_n500_n697# a_n558_n600# w_n758_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=5
C0 w_n758_n897# a_n558_n600# 0.361528f
C1 w_n758_n897# a_n500_n697# 1.61638f
C2 a_500_n600# w_n758_n897# 0.361528f
C3 a_n558_n600# a_n500_n697# 0.243898f
C4 a_500_n600# a_n558_n600# 0.079546f
C5 a_500_n600# a_n500_n697# 0.243898f
C6 a_500_n600# 0 0.402067f
C7 a_n558_n600# 0 0.402067f
C8 a_n500_n697# 0 1.41779f
C9 w_n758_n897# 0 9.64891f
.ends

.subckt trans_gate in ena_b ena out avdd vss
XXM1 ena out vss in sky130_fd_pr__nfet_g5v0d10v5_69BJMM
XXM2 avdd out ena_b in vss sky130_fd_pr__pfet_g5v0d10v5_E7V9VM
C0 ena_b ena 0.040022f
C1 ena out 0.455968f
C2 ena_b in 0.484944f
C3 ena_b avdd 0.458648f
C4 out in 0.395476f
C5 avdd out 0.18948f
C6 ena_b out 0.781385f
C7 ena in 0.435683f
C8 avdd ena 0.062182f
C9 avdd in 0.273851f
C10 in vss 0.96413f
C11 out vss 1.721452f
C12 ena_b vss 1.715065f
C13 avdd vss 9.963131f
C14 ena vss 3.308732f
.ends

.subckt sky130_fd_pr__pfet_01v8_C2YSV5 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
+ 0
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
C0 a_n300_n197# w_n496_n319# 1.05203f
C1 a_n358_n100# a_n300_n197# 0.042408f
C2 a_n300_n197# a_300_n100# 0.042408f
C3 a_n358_n100# w_n496_n319# 0.085201f
C4 a_300_n100# w_n496_n319# 0.085201f
C5 a_n358_n100# a_300_n100# 0.021684f
C6 a_300_n100# 0 0.071857f
C7 a_n358_n100# 0 0.071857f
C8 a_n300_n197# 0 0.838987f
C9 w_n496_n319# 0 2.60523f
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9E5 w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
+ 0
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n100_n197# w_n296_n319# 0.434431f
C1 a_n158_n100# a_n100_n197# 0.026809f
C2 a_n100_n197# a_100_n100# 0.026809f
C3 a_n158_n100# w_n296_n319# 0.085221f
C4 a_100_n100# w_n296_n319# 0.085221f
C5 a_n158_n100# a_100_n100# 0.055609f
C6 a_100_n100# 0 0.060699f
C7 a_n158_n100# 0 0.060699f
C8 a_n100_n197# 0 0.310981f
C9 w_n296_n319# 0 1.64714f
.ends

.subckt sky130_fd_pr__pfet_01v8_GGMWVD w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
+ 0
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
C0 a_n800_n197# w_n996_n319# 2.59374f
C1 a_n858_n100# a_n800_n197# 0.049339f
C2 a_n800_n197# a_800_n100# 0.049339f
C3 a_n858_n100# w_n996_n319# 0.085193f
C4 a_800_n100# w_n996_n319# 0.085193f
C5 a_800_n100# 0 0.091337f
C6 a_n858_n100# 0 0.091337f
C7 a_n800_n197# 0 2.159f
C8 w_n996_n319# 0 5.00228f
.ends

.subckt sky130_fd_pr__pfet_01v8_CDT3CS a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
+ 0
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
C0 a_n1600_n197# w_n1796_n319# 5.05964f
C1 a_n1658_n100# a_n1600_n197# 0.049339f
C2 a_n1600_n197# a_1600_n100# 0.049339f
C3 a_n1658_n100# w_n1796_n319# 0.085193f
C4 a_1600_n100# w_n1796_n319# 0.085193f
C5 a_1600_n100# 0 0.091337f
C6 a_n1658_n100# 0 0.091337f
C7 a_n1600_n197# 0 4.27103f
C8 w_n1796_n319# 0 8.81803f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
C0 a_n158_n100# a_n100_n188# 0.026809f
C1 a_100_n100# a_n158_n100# 0.055609f
C2 a_100_n100# a_n100_n188# 0.026809f
C3 a_100_n100# a_n292_n322# 0.137447f
C4 a_n158_n100# a_n292_n322# 0.137447f
C5 a_n100_n188# a_n292_n322# 0.688242f
.ends

.subckt sky130_fd_pr__pfet_01v8_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397# a_100_n300#
+ 0
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
C0 a_n100_n397# w_n296_n519# 0.434431f
C1 a_n158_n300# a_n100_n397# 0.069551f
C2 a_n100_n397# a_100_n300# 0.069551f
C3 a_n158_n300# w_n296_n519# 0.207171f
C4 a_100_n300# w_n296_n519# 0.207171f
C5 a_n158_n300# a_100_n300# 0.164742f
C6 a_100_n300# 0 0.161554f
C7 a_n158_n300# 0 0.161554f
C8 a_n100_n397# 0 0.328882f
C9 w_n296_n519# 0 2.55335f
.ends

.subckt sky130_fd_pr__nfet_01v8_697RXD a_800_n100# a_n858_n100# a_n800_n188# a_n960_n274#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n960_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
C0 a_n858_n100# a_n800_n188# 0.049339f
C1 a_800_n100# a_n800_n188# 0.049339f
C2 a_800_n100# a_n960_n274# 0.176968f
C3 a_n858_n100# a_n960_n274# 0.176968f
C4 a_n800_n188# a_n960_n274# 4.65384f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_4T6WVE a_100_n130# a_n292_n352# a_n158_n130#
+ a_n100_n218#
X0 a_100_n130# a_n100_n218# a_n158_n130# a_n292_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=1
C0 a_n158_n130# a_n100_n218# 0.033221f
C1 a_100_n130# a_n158_n130# 0.071979f
C2 a_100_n130# a_n100_n218# 0.033221f
C3 a_100_n130# a_n292_n352# 0.168646f
C4 a_n158_n130# a_n292_n352# 0.168646f
C5 a_n100_n218# a_n292_n352# 0.692382f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_6975WM a_800_n130# a_n992_n352# a_n858_n130#
+ a_n800_n218#
X0 a_800_n130# a_n800_n218# a_n858_n130# a_n992_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
C0 a_n858_n130# a_n800_n218# 0.061878f
C1 a_800_n130# a_n800_n218# 0.061878f
C2 a_800_n130# a_n992_n352# 0.209212f
C3 a_n858_n130# a_n992_n352# 0.209212f
C4 a_n800_n218# a_n992_n352# 4.43441f
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DEN7YK a_800_n100# a_n992_n322# a_n858_n100#
+ a_n800_n188#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n992_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
C0 a_n858_n100# a_n800_n188# 0.049339f
C1 a_800_n100# a_n800_n188# 0.049339f
C2 a_800_n100# a_n992_n322# 0.168056f
C3 a_n858_n100# a_n992_n322# 0.168056f
C4 a_n800_n188# a_n992_n322# 4.39578f
.ends

.subckt sky130_fd_pr__pfet_01v8_G3L97A w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
+ 0
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
C0 a_n800_n197# w_n996_n319# 2.59374f
C1 a_n858_n100# a_n800_n197# 0.049339f
C2 a_n800_n197# a_800_n100# 0.049339f
C3 a_n858_n100# w_n996_n319# 0.085193f
C4 a_800_n100# w_n996_n319# 0.085193f
C5 a_800_n100# 0 0.091337f
C6 a_n858_n100# 0 0.091337f
C7 a_n800_n197# 0 2.159f
C8 w_n996_n319# 0 5.00228f
.ends

.subckt sky130_fd_pr__nfet_01v8_C8TQ3N a_n158_n300# a_n100_n388# a_n260_n474# a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n260_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
C0 a_n158_n300# a_n100_n388# 0.069551f
C1 a_100_n300# a_n158_n300# 0.164742f
C2 a_100_n300# a_n100_n388# 0.069551f
C3 a_100_n300# a_n260_n474# 0.369164f
C4 a_n158_n300# a_n260_n474# 0.369164f
C5 a_n100_n388# a_n260_n474# 0.742994f
.ends

.subckt comp_hyst vref ibias net2 ena net5 vin dvss net1 ena_b dvdd out net3 net4
XXMD16[0] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXM12 dvss net1 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
XXM14 dvss net2 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXM13 dvss net5 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
Xx1 ibias ena_b ena net5 dvdd dvss trans_gate
XXM15 ena net4 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_C2YSV5
XXM16 ena net3 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_C2YSV5
XXM17 dvss out ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXMD1[19] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM18 ena ena_b dvdd dvdd dvss sky130_fd_pr__pfet_01v8_C2YSV5
XXMD1[18] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM19 dvss ena_b ena dvss sky130_fd_pr__nfet_01v8_V433WY
XXM6[3] net3 net4 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXM3[1] dvdd net4 net4 dvdd dvss sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[17] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[2] net3 net4 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_CDT3CS
XXM3[0] dvdd net4 net4 dvdd dvss sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[16] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[1] net3 net4 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXM6[0] net3 net4 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_CDT3CS
XXMD1[15] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[13] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[14] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[9] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[12] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[8] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[11] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[7] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[10] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[6] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[4] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[5] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XD1 dvss vref sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[3] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM7 dvdd net4 net2 dvdd dvss sky130_fd_pr__pfet_01v8_GGMWVD
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[2] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM9 dvdd dvdd net3 out dvss sky130_fd_pr__pfet_01v8_3HBZVM
XXM8 dvss net2 net2 dvss sky130_fd_pr__nfet_01v8_697RXD
XXMDN13[7] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXM1[1] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXMD1[1] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM1[0] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM4[1] net3 net3 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXMDN13[6] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMD1[0] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_J2L9E5
XXM4[0] net3 net3 dvdd dvdd dvss sky130_fd_pr__pfet_01v8_CDT3CS
XXMDN13[5] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[4] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN8[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMDN8[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMD16[5] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXMD16[4] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[1] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[1] dvdd net4 net3 dvdd dvss sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[3] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[0] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[0] dvdd net4 net3 dvdd dvss sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[2] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXMD8[1] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_G3L97A
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 dvss vin sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXM10 out net2 dvss dvss sky130_fd_pr__nfet_01v8_C8TQ3N
XXMD8[0] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_G3L97A
XXMD16[1] dvdd dvdd dvdd dvdd dvss sky130_fd_pr__pfet_01v8_XTWSDC
XXM11 dvss net5 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
C0 out net2 1.07639f
C1 vref net4 1.76685f
C2 ena ibias 0.077568f
C3 net2 net5 0.140511f
C4 ena_b ibias 0.081201f
C5 vin vref 1.678694f
C6 net2 net4 1.045614f
C7 out net5 0.038132f
C8 net1 net5 2.752974f
C9 dvdd ibias 0.013497f
C10 vref net3 1.084347f
C11 net2 ena 0.032097f
C12 out net4 0.385987f
C13 net2 ena_b 0.527846f
C14 net1 net4 0.063495f
C15 net4 net5 0.078978f
C16 net2 net3 0.354659f
C17 vin net1 0.622826f
C18 ena net1 0.02159f
C19 out ena_b 0.483538f
C20 ena net5 1.030568f
C21 dvdd net2 0.465128f
C22 ena_b net5 1.036401f
C23 vin net4 0.071217f
C24 out net3 1.498908f
C25 net3 net5 0.010117f
C26 ena net4 0.798922f
C27 ena_b net4 0.014856f
C28 net4 net3 17.40976f
C29 out dvdd 0.989102f
C30 dvdd net5 0.064156f
C31 vin net3 0.502438f
C32 ena_b ena 2.479058f
C33 dvdd net4 16.580809f
C34 ena net3 0.467559f
C35 ena_b net3 0.012875f
C36 ibias net5 0.083723f
C37 dvdd ena 2.004081f
C38 dvdd ena_b 0.515966f
C39 vref net1 1.239698f
C40 dvdd net3 14.160767f
C41 vref net5 0.019445f
C42 net3 dvss 21.002346f
C43 vin dvss 9.844718f
C44 net1 dvss 4.887807f
C45 net4 dvss 11.991661f
C46 vref dvss 10.502412f
C47 out dvss 3.311475f
C48 ibias dvss 0.799971f
C49 net5 dvss 26.223053f
C50 ena_b dvss 9.433245f
C51 dvdd dvss 0.179918p
C52 ena dvss 7.901359f
C53 net2 dvss 7.398622f
.ends

.subckt sky130_vbl_ip__overvoltage avdd dvdd ena vtrip[3] ibias vtrip[2] ovout vbg
+ vtrip[1] vtrip[0] dvss avss
Xvoltage_divider_0 multiplexer_0/in_0000 multiplexer_0/in_0001 multiplexer_0/in_0010
+ multiplexer_0/in_0011 multiplexer_0/in_0101 multiplexer_0/in_0110 multiplexer_0/in_0111
+ multiplexer_0/in_1001 multiplexer_0/in_1010 multiplexer_0/in_1011 multiplexer_0/in_1101
+ multiplexer_0/in_1111 ena voltage_divider_0/m1_7155_3601# voltage_divider_0/m1_10901_8137#
+ voltage_divider_0/m1_7155_14563# voltage_divider_0/m1_7691_16075# voltage_divider_0/m1_3399_9649#
+ voltage_divider_0/m1_10911_2089# voltage_divider_0/m1_7155_3223# voltage_divider_0/m1_3399_12673#
+ voltage_divider_0/m1_10911_15697# voltage_divider_0/m1_3399_3979# voltage_divider_0/m1_7155_5491#
+ voltage_divider_0/m1_3399_7381# voltage_divider_0/m1_7155_9271# voltage_divider_0/m1_10911_13429#
+ voltage_divider_0/m1_7155_12295# voltage_divider_0/m1_7691_14563# voltage_divider_0/m1_3399_16453#
+ voltage_divider_0/m1_7155_7759# voltage_divider_0/m1_3935_10405# voltage_divider_0/m1_179_3979#
+ voltage_divider_0/51 voltage_divider_0/m1_7155_10027# voltage_divider_0/m1_3399_199#
+ voltage_divider_0/m1_3399_3601# voltage_divider_0/m1_179_13051# voltage_divider_0/m1_3935_14185#
+ voltage_divider_0/m1_179_199# voltage_divider_0/m1_7691_9271# voltage_divider_0/m1_7691_12295#
+ voltage_divider_0/m1_7155_10783# voltage_divider_0/m1_3935_4357# voltage_divider_0/m1_7691_10027#
+ voltage_divider_0/m1_7155_7003# voltage_divider_0/m1_3399_15697# voltage_divider_0/m1_3935_8137#
+ voltage_divider_0/m1_3399_955# voltage_divider_0/m1_7691_10783# voltage_divider_0/m1_179_12295#
+ voltage_divider_0/m1_7155_16831# voltage_divider_0/m1_179_955# voltage_divider_0/m1_7691_7003#
+ voltage_divider_0/m1_179_6247# voltage_divider_0/m1_7155_955# voltage_divider_0/m1_3399_2467#
+ voltage_divider_0/m1_179_16075# voltage_divider_0/m1_3935_8893# voltage_divider_0/m1_3935_11917#
+ voltage_divider_0/m1_179_2467# voltage_divider_0/m1_3935_5113# voltage_divider_0/m1_7155_2845#
+ voltage_divider_0/m1_10911_16453# voltage_divider_0/m1_3399_13429# voltage_divider_0/m1_7155_13051#
+ voltage_divider_0/m1_10911_1333# voltage_divider_0/m1_179_16831# voltage_divider_0/m1_179_10027#
+ voltage_divider_0/m1_7155_4735# voltage_divider_0/m1_3399_17209# voltage_divider_0/m1_10911_14185#
+ voltage_divider_0/m1_179_7003# voltage_divider_0/m1_3399_3223# voltage_divider_0/m1_3399_6625#
+ voltage_divider_0/m1_3935_9649# voltage_divider_0/m1_10911_11917# voltage_divider_0/m1_7691_13051#
+ voltage_divider_0/m1_179_3223# voltage_divider_0/m1_3935_12673# voltage_divider_0/m1_3399_2845#
+ multiplexer_0/in_1100 voltage_divider_0/m1_10911_12673# voltage_divider_0/m1_3935_7381#
+ voltage_divider_0/m1_3935_16453# avdd voltage_divider_0/m1_7155_577# voltage_divider_0/m1_7155_17209#
+ voltage_divider_0/m1_3399_5869# voltage_divider_0/m1_179_10783# voltage_divider_0/m1_7155_199#
+ voltage_divider_0/m1_3399_11161# voltage_divider_0/m1_3399_14941# voltage_divider_0/m1_3399_2089#
+ voltage_divider_0/m1_7155_2467# voltage_divider_0/m1_179_14563# voltage_divider_0/m1_7155_8515#
+ voltage_divider_0/m1_7155_15319# voltage_divider_0/m1_3935_15697# voltage_divider_0/m1_179_5491#
+ voltage_divider_0/m1_3399_1711# voltage_divider_0/m1_7155_2089# voltage_divider_0/m1_179_1711#
+ multiplexer_0/in_0100 voltage_divider_0/m1_7691_15319# voltage_divider_0/m1_3399_10405#
+ voltage_divider_0/m1_179_13807# voltage_divider_0/m1_7155_3979# voltage_divider_0/m1_7155_13807#
+ voltage_divider_0/m1_3399_14185# voltage_divider_0/m1_7155_6247# voltage_divider_0/m1_10911_2845#
+ voltage_divider_0/m1_7155_11539# voltage_divider_0/m1_179_9271# voltage_divider_0/m1_3399_4357#
+ voltage_divider_0/m1_3935_13429# multiplexer_0/in_1110 voltage_divider_0/m1_7691_13807#
+ voltage_divider_0/m1_179_7759# voltage_divider_0/m1_3399_577# voltage_divider_0/m1_3399_8137#
+ multiplexer_0/in_1000 voltage_divider_0/m1_3935_6625# voltage_divider_0/m1_3399_8893#
+ voltage_divider_0/m1_179_11539# voltage_divider_0/m1_3399_11917# voltage_divider_0/m1_3399_5113#
+ voltage_divider_0/m1_179_15319# voltage_divider_0/m1_10911_577# voltage_divider_0/m1_7155_1711#
+ voltage_divider_0/m1_7155_16075# voltage_divider_0/m1_3399_1333# voltage_divider_0/m1_3935_5869#
+ voltage_divider_0/m1_10911_14941# voltage_divider_0/m1_10901_199# voltage_divider_0/m1_7155_1333#
+ voltage_divider_0/m1_179_4735# voltage_divider_0/m1_179_8515# voltage_divider_0/m1_3935_11161#
+ voltage_divider_0/m1_3935_14941# avss voltage_divider
Xmultiplexer_0 multiplexer_0/in_0000 multiplexer_0/in_0001 multiplexer_0/in_0011 multiplexer_0/in_0100
+ multiplexer_0/in_0101 multiplexer_0/in_0110 level_shifter_3/out level_shifter_3/out_b
+ level_shifter_2/out vin level_shifter_1/out_b multiplexer_0/in_1000 multiplexer_0/in_1001
+ multiplexer_0/in_1010 multiplexer_0/in_1100 multiplexer_0/in_1101 multiplexer_0/in_1110
+ multiplexer_0/in_1111 multiplexer_0/trans_gate_m_37/in multiplexer_0/trans_gate_m_32/in
+ level_shifter_0/out_b multiplexer_0/trans_gate_m_7/out multiplexer_0/in_1011 multiplexer_0/trans_gate_m_27/in
+ multiplexer_0/trans_gate_m_3/out multiplexer_0/trans_gate_m_33/in multiplexer_0/trans_gate_m_34/in
+ multiplexer_0/trans_gate_m_28/in multiplexer_0/in_0111 multiplexer_0/in_0010 multiplexer_0/trans_gate_m_5/out
+ multiplexer_0/trans_gate_m_20/in multiplexer_0/trans_gate_m_31/in multiplexer_0/trans_gate_m_23/in
+ multiplexer_0/trans_gate_m_9/out level_shifter_2/out_b multiplexer_0/trans_gate_m_29/in
+ avss level_shifter_1/out level_shifter_0/out avdd multiplexer
Xlevel_shifter_0 vtrip[0] level_shifter_0/out level_shifter_0/out_b dvss level_shifter_0/in_b
+ avss dvdd avdd level_shifter
Xlevel_shifter_1 vtrip[1] level_shifter_1/out level_shifter_1/out_b dvss level_shifter_1/in_b
+ avss dvdd avdd level_shifter
Xlevel_shifter_2 vtrip[2] level_shifter_2/out level_shifter_2/out_b dvss level_shifter_2/in_b
+ avss dvdd avdd level_shifter
Xlevel_shifter_3 vtrip[3] level_shifter_3/out level_shifter_3/out_b dvss level_shifter_3/in_b
+ avss dvdd avdd level_shifter
Xcomp_hyst_0 vbg ibias comp_hyst_0/net2 ena comp_hyst_0/net5 vin dvss comp_hyst_0/net1
+ comp_hyst_0/ena_b dvdd ovout comp_hyst_0/net3 comp_hyst_0/net4 comp_hyst
C1 vin level_shifter_0/out_b 0.104612f
C2 multiplexer_0/in_0011 avdd 0.020365f
C3 vtrip[2] avdd 0.182561f
C4 level_shifter_1/out_b level_shifter_2/out_b 0.42065f
C5 level_shifter_3/out_b avdd 0.152807f
C6 level_shifter_2/out_b avss 4.656484f
C7 ena level_shifter_2/in_b 0.018249f
C8 level_shifter_2/out avdd 0.917194f
C9 initials_0/m4_3195_879# initials_0/m4_2307_879# 0.186835f
C10 avss multiplexer_0/trans_gate_m_34/in 1.015015f
C11 level_shifter_1/out multiplexer_0/trans_gate_m_27/in 0.150564f
C12 level_shifter_0/out_b multiplexer_0/trans_gate_m_33/in 0.191061f
C13 multiplexer_0/in_1011 multiplexer_0/in_1110 0.062764f
C14 voltage_divider_0/m1_7155_199# avss 0.079556f
C15 multiplexer_0/in_0001 multiplexer_0/in_0000 0.694704f
C16 avss voltage_divider_0/m1_7155_3223# 0.079556f
C17 level_shifter_2/in_b avdd 0.084148f
C18 voltage_divider_0/m1_3399_6625# avss 0.092648f
C19 dvdd level_shifter_0/in_b 0.583879f
C20 voltage_divider_0/m1_3399_12673# avss 0.092648f
C21 vtrip[0] dvdd 3.623714f
C22 avss multiplexer_0/trans_gate_m_9/out 0.824159f
C23 multiplexer_0/in_0110 multiplexer_0/in_1000 0.013534f
C24 level_shifter_3/in_b vtrip[1] 0.112568f
C25 avss dvdd 0.303163f
C26 avdd multiplexer_0/in_1010 0.102314f
C27 avss voltage_divider_0/m1_10911_12673# 0.092648f
C28 avss voltage_divider_0/m1_10901_8137# 0.096787f
C29 level_shifter_0/out multiplexer_0/in_0011 0.022222f
C30 vin initials_0/m4_2474_2379# 0.030085f
C31 initials_0/m4_2374_1229# initials_0/m4_2307_879# 0.249242f
C32 avss multiplexer_0/in_1101 1.332217f
C33 level_shifter_0/out level_shifter_2/out 0.116748f
C34 ovout dvdd 0.172896f
C35 comp_hyst_0/net4 dvdd 0.014075f
C36 ena vtrip[1] 0.370865f
C37 multiplexer_0/in_0100 avss 1.737438f
C39 avss voltage_divider_0/m1_3399_14185# 0.092648f
C40 avss voltage_divider_0/m1_10911_1333# 0.092648f
C41 multiplexer_0/in_0000 multiplexer_0/in_0010 0.704f
C42 voltage_divider_0/m1_10911_14185# avss 0.092648f
C43 level_shifter_3/in_b ena 0.018249f
C44 multiplexer_0/in_1000 avdd 0.243334f
C45 initials_0/m4_1419_2382# initials_0/m4_1419_879# 0.012147f
C46 avss voltage_divider_0/m1_7155_13807# 0.092648f
C47 vtrip[1] avdd 0.139709f
C48 multiplexer_0/in_0001 multiplexer_0/in_0011 0.550521f
C49 level_shifter_1/out avdd 1.674446f
C50 avss voltage_divider_0/m1_3399_3979# 0.094199f
C51 voltage_divider_0/m1_3399_9649# avss 0.092648f
C52 avss voltage_divider_0/m1_7155_10027# 0.092648f
C53 voltage_divider_0/m1_10911_14941# avss 0.092648f
C54 multiplexer_0/in_0101 multiplexer_0/in_1010 0.017461f
C55 level_shifter_3/in_b avdd 0.083435f
C56 avss voltage_divider_0/m1_179_7003# 0.092648f
C57 multiplexer_0/in_0110 avdd 0.017654f
C58 avss multiplexer_0/trans_gate_m_31/in 0.842496f
C59 avss multiplexer_0/trans_gate_m_7/out 0.685192f
C60 multiplexer_0/trans_gate_m_28/in level_shifter_1/out_b 0.229406f
C61 avss voltage_divider_0/m1_179_15319# 0.092648f
C62 multiplexer_0/trans_gate_m_28/in avss 0.591114f
C63 voltage_divider_0/m1_3935_8137# avss 0.092648f
C64 level_shifter_0/out multiplexer_0/trans_gate_m_29/in 0.039227f
C65 multiplexer_0/trans_gate_m_23/in multiplexer_0/in_1010 0.025395f
C66 voltage_divider_0/m1_7155_5491# avss 0.091766f
C67 initials_0/m4_1419_879# initials_0/m4_2307_879# 0.186835f
C68 level_shifter_0/out multiplexer_0/trans_gate_m_27/in 0.01968f
C69 vtrip[0] level_shifter_0/in_b 0.084412f
C70 voltage_divider_0/m1_179_955# avss 0.092648f
C71 avss level_shifter_0/in_b 0.797957f
C72 ena avdd 0.103523f
C73 avss vtrip[0] 0.836718f
C74 level_shifter_1/out_b avss 6.407568f
C75 vin dvdd 1.159184f
C76 voltage_divider_0/m1_7155_2845# avss 0.079556f
C77 avss multiplexer_0/in_1001 0.630282f
C78 multiplexer_0/in_0011 multiplexer_0/in_0010 1.712367f
C79 vin comp_hyst_0/net5 0.017967f
C80 avss voltage_divider_0/m1_7155_16075# 0.092648f
C81 multiplexer_0/in_0101 multiplexer_0/in_1000 0.210796f
C82 ibias dvdd 4.225524f
C83 voltage_divider_0/m1_7691_12295# avss 0.092648f
C84 level_shifter_0/out level_shifter_1/out 0.728282f
C85 initials_0/m4_2374_1229# initials_0/m4_1419_1229# 0.119924f
C86 ibias comp_hyst_0/net5 0.148155f
C87 avss voltage_divider_0/m1_7155_8515# 0.091766f
C88 voltage_divider_0/m1_179_7759# avss 0.092648f
C89 voltage_divider_0/m1_179_11539# avss 0.092648f
C90 voltage_divider_0/m1_10911_13429# avss 0.092648f
C91 vtrip[2] vtrip[3] 2.127573f
C92 multiplexer_0/in_1011 avss 0.726547f
C93 multiplexer_0/in_0110 multiplexer_0/in_0101 0.412123f
C94 avss voltage_divider_0/m1_3935_15697# 0.092648f
C95 multiplexer_0/in_1011 multiplexer_0/in_1001 0.302679f
C96 level_shifter_0/out_b level_shifter_2/out 0.126128f
C97 avss voltage_divider_0/m1_3399_199# 0.079556f
C100 voltage_divider_0/m1_10911_2845# avss 0.092648f
C101 level_shifter_2/in_b vtrip[3] 0.087257f
C102 multiplexer_0/trans_gate_m_20/in avss 0.769866f
C103 voltage_divider_0/m1_3399_5113# avss 0.092648f
C104 voltage_divider_0/m1_10911_577# avss 0.092648f
C105 avss voltage_divider_0/m1_3399_11161# 0.092648f
C106 voltage_divider_0/m1_179_6247# avss 0.092648f
C107 level_shifter_3/out level_shifter_3/out_b 0.706827f
C108 level_shifter_3/out level_shifter_2/out 0.203516f
C109 level_shifter_0/out avdd 1.59437f
C110 voltage_divider_0/m1_3935_11161# avss 0.092648f
C111 avss voltage_divider_0/m1_3399_11917# 0.092648f
C112 multiplexer_0/in_0101 avdd 0.150109f
C113 voltage_divider_0/m1_179_3979# avss 0.092648f
C114 avss voltage_divider_0/m1_3935_5869# 0.092648f
C115 level_shifter_0/out_b multiplexer_0/in_1010 0.052242f
C116 initials_0/m4_1419_879# initials_0/m4_1419_1229# 0.213636f
C117 vin level_shifter_0/in_b 0.174826f
C118 vin vtrip[0] 0.335778f
C119 vin level_shifter_1/out_b 0.286622f
C120 vin avss 2.130694f
C121 voltage_divider_0/m1_179_3223# avss 0.092648f
C122 avss voltage_divider_0/m1_3399_955# 0.079556f
C123 ibias level_shifter_0/in_b 0.079403f
C124 voltage_divider_0/51 avss 0.092648f
C125 ibias vtrip[0] 0.098883f
C126 avss ibias 0.011481f
C127 voltage_divider_0/m1_3935_5113# avss 0.092648f
C128 level_shifter_1/out_b multiplexer_0/trans_gate_m_33/in 0.240574f
C129 level_shifter_0/out_b multiplexer_0/trans_gate_m_27/in 0.184967f
C130 multiplexer_0/trans_gate_m_33/in avss 1.158379f
C131 avss voltage_divider_0/m1_3399_5869# 0.092648f
C132 initials_0/m4_2474_2379# initials_0/m4_2374_1229# 0.213636f
C133 voltage_divider_0/m1_3935_16453# avss 0.092648f
C134 multiplexer_0/in_0001 avdd 0.087327f
C135 vtrip[1] vtrip[3] 0.374288f
C136 voltage_divider_0/m1_3399_10405# avss 0.092648f
C137 comp_hyst_0/net4 ibias 0.049422f
C138 avss voltage_divider_0/m1_3935_14941# 0.092648f
C139 level_shifter_0/out_b level_shifter_1/out 1.909585f
C140 multiplexer_0/in_0000 multiplexer_0/in_0100 0.028175f
C141 initials_0/m4_2474_2379# initials_0/m4_3195_2379# 0.248819f
C142 level_shifter_3/in_b vtrip[3] 0.214591f
C143 level_shifter_3/out_b level_shifter_2/out_b 0.322285f
C144 avss voltage_divider_0/m1_3399_16453# 0.092648f
C146 level_shifter_2/out_b level_shifter_2/out 0.729726f
C147 avss voltage_divider_0/m1_3935_10405# 0.092648f
C148 avss voltage_divider_0/m1_3935_11917# 0.092648f
C149 multiplexer_0/in_0110 level_shifter_0/out_b 0.200806f
C150 multiplexer_0/in_1111 avdd 0.012402f
C151 level_shifter_3/out_b multiplexer_0/trans_gate_m_34/in 0.245053f
C152 avss voltage_divider_0/m1_179_13051# 0.092648f
C153 level_shifter_2/out multiplexer_0/trans_gate_m_34/in 0.19431f
C154 multiplexer_0/in_0111 multiplexer_0/in_1010 0.78608f
C155 avss voltage_divider_0/m1_7691_10783# 0.092648f
C156 avss voltage_divider_0/m1_3935_7381# 0.092648f
C157 multiplexer_0/in_1110 multiplexer_0/in_1010 0.01934f
C158 level_shifter_1/in_b dvdd 0.574098f
C159 ena vtrip[3] 0.396701f
C160 avdd multiplexer_0/in_0010 0.026116f
C161 initials_0/m4_1419_2382# initials_0/m4_1419_1229# 0.099027f
C162 vtrip[2] dvdd 1.88741f
C163 voltage_divider_0/m1_10911_16453# avss 0.091285f
C164 initials_0/m4_3395_1229# initials_0/m4_3195_879# 0.122517f
C165 avdd vtrip[3] 0.301175f
C166 level_shifter_0/out_b avdd 1.528315f
C167 avss voltage_divider_0/m1_7155_1333# 0.079556f
C168 avss voltage_divider_0/m1_3399_2845# 0.079556f
C169 dvdd comp_hyst_0/net3 0.053947f
C170 vin ibias 0.021594f
C171 multiplexer_0/in_0111 multiplexer_0/in_1000 0.303441f
C172 multiplexer_0/in_0000 avss 2.026233f
C173 multiplexer_0/in_0100 multiplexer_0/in_0011 0.172839f
C174 avss voltage_divider_0/m1_10911_2089# 0.092648f
C175 avss voltage_divider_0/m1_3935_12673# 0.092648f
C176 dvdd level_shifter_2/in_b 0.573131f
C177 avss voltage_divider_0/m1_179_12295# 0.092648f
C178 voltage_divider_0/m1_10911_15697# avss 0.092648f
C179 avss voltage_divider_0/m1_3399_13429# 0.092648f
C180 multiplexer_0/in_0110 multiplexer_0/in_0111 1.257687f
C181 level_shifter_3/out avdd 0.328925f
C182 level_shifter_1/out level_shifter_2/out_b 0.13455f
C183 avss voltage_divider_0/m1_7155_955# 0.079556f
C184 voltage_divider_0/m1_7155_15319# avss 0.092648f
C185 initials_0/m4_2374_1229# initials_0/m4_3395_1229# 0.216092f
C186 voltage_divider_0/m1_7155_7003# avss 0.092648f
C187 avss voltage_divider_0/m1_3399_14941# 0.092648f
C188 voltage_divider_0/m1_3935_4357# avss 0.092648f
C189 level_shifter_1/in_b vtrip[0] 0.151155f
C190 voltage_divider_0/m1_3399_1711# avss 0.079556f
C191 avss voltage_divider_0/m1_7155_7759# 0.091766f
C192 level_shifter_0/out level_shifter_0/out_b 1.951787f
C193 level_shifter_1/in_b avss 1.062538f
C194 avss voltage_divider_0/m1_179_199# 0.092648f
C195 initials_0/m4_1419_2382# initials_0/m4_2474_2379# 0.449761f
C196 multiplexer_0/in_0001 multiplexer_0/in_0010 0.278453f
C197 multiplexer_0/in_0111 avdd 0.063929f
C198 avss multiplexer_0/in_0011 1.019819f
C199 initials_0/m4_3395_1229# initials_0/m4_3195_2379# 0.213636f
C200 multiplexer_0/in_1110 avdd 0.010472f
C201 vtrip[2] vtrip[0] 0.582856f
C202 vtrip[2] avss 1.340418f
C203 dvdd vtrip[1] 2.077883f
C204 level_shifter_1/out_b level_shifter_3/out_b 0.033854f
C205 level_shifter_3/out_b avss 3.685153f
C206 level_shifter_1/out_b level_shifter_2/out 0.195073f
C207 avss level_shifter_2/out 4.962986f
C208 voltage_divider_0/m1_3399_3223# avss 0.079556f
C209 level_shifter_3/in_b dvdd 0.066238f
C210 voltage_divider_0/m1_179_16075# avss 0.092648f
C211 voltage_divider_0/m1_7155_1711# avss 0.079556f
C212 level_shifter_2/out_b avdd 0.598585f
C213 vtrip[0] level_shifter_2/in_b 0.119187f
C214 avss level_shifter_2/in_b 1.063496f
C215 voltage_divider_0/m1_7155_2089# avss 0.079556f
C216 ena dvdd 0.178439f
C217 avss multiplexer_0/in_1010 0.960204f
C218 multiplexer_0/in_0110 multiplexer_0/in_0100 0.622562f
C219 level_shifter_0/out_b multiplexer_0/trans_gate_m_3/out 0.314969f
C220 avss voltage_divider_0/m1_3399_2089# 0.079556f
C221 multiplexer_0/in_1010 multiplexer_0/in_1001 0.528857f
C222 voltage_divider_0/m1_7155_2467# avss 0.079556f
C223 vbg dvdd 0.107944f
C224 level_shifter_0/out multiplexer_0/in_0111 0.038449f
C225 multiplexer_0/in_0111 multiplexer_0/in_0101 0.47148f
C226 avss multiplexer_0/trans_gate_m_37/in 0.899199f
C227 voltage_divider_0/m1_3399_8893# avss 0.092648f
C228 dvdd avdd 0.213897f
C229 avss multiplexer_0/trans_gate_m_29/in 0.673122f
C230 avss multiplexer_0/trans_gate_m_27/in 0.854834f
C231 level_shifter_0/out_b multiplexer_0/in_0010 0.010603f
C232 dvdd rocket_0/m1_n9_n9# 0.089427f
C233 multiplexer_0/trans_gate_m_28/in level_shifter_1/out 0.459668f
C234 level_shifter_0/out level_shifter_2/out_b 0.406705f
C235 multiplexer_0/in_1011 multiplexer_0/in_1010 0.845489f
C236 voltage_divider_0/m1_3935_13429# avss 0.092648f
C237 avdd multiplexer_0/in_1101 0.068496f
C238 voltage_divider_0/m1_179_10027# avss 0.092648f
C239 voltage_divider_0/m1_7155_4735# avss 0.091766f
C240 avss voltage_divider_0/m1_7691_13051# 0.092648f
C241 avss multiplexer_0/in_1000 1.337429f
C242 level_shifter_0/in_b vtrip[1] 0.012661f
C243 vtrip[0] vtrip[1] 3.223579f
C244 multiplexer_0/in_1000 multiplexer_0/in_1001 0.476548f
C245 multiplexer_0/in_0100 avdd 0.113418f
C246 avss vtrip[1] 1.234469f
C247 level_shifter_1/out_b level_shifter_1/out 2.402098f
C248 level_shifter_1/out avss 7.17497f
C249 multiplexer_0/in_1110 multiplexer_0/in_1100 0.235044f
C250 voltage_divider_0/m1_179_1711# avss 0.092648f
C251 level_shifter_3/in_b vtrip[0] 0.121954f
C252 avss voltage_divider_0/m1_3399_2467# 0.079556f
C253 level_shifter_3/in_b avss 1.099654f
C254 voltage_divider_0/m1_179_2467# avss 0.092648f
C255 voltage_divider_0/m1_7155_577# avss 0.079556f
C256 multiplexer_0/in_0110 avss 0.953726f
C257 level_shifter_0/out dvdd 0.110033f
C258 voltage_divider_0/m1_7691_14563# avss 0.092648f
C259 ibias comp_hyst_0/net3 0.176846f
C260 multiplexer_0/in_1011 multiplexer_0/in_1000 0.026096f
C261 multiplexer_0/in_1111 multiplexer_0/in_1110 0.084259f
C262 vtrip[0] ena 0.314015f
C263 vin initials_0/m4_3195_2379# 0.043283f
C264 avss ena 6.551044f
C265 voltage_divider_0/m1_10911_11917# avss 0.092648f
C266 avss voltage_divider_0/m1_3935_9649# 0.092648f
C268 voltage_divider_0/m1_7691_15319# avss 0.092648f
C269 voltage_divider_0/m1_7691_7003# avss 0.092648f
C270 avss voltage_divider_0/m1_7691_9271# 0.092648f
C271 multiplexer_0/in_0101 multiplexer_0/in_0100 0.508949f
C272 level_shifter_0/in_b avdd 0.094194f
C273 vtrip[0] avdd 0.184643f
C274 level_shifter_1/out_b avdd 1.053612f
C275 avss voltage_divider_0/m1_7155_3979# 0.091766f
C276 avss avdd 1.608667p
C277 avdd multiplexer_0/in_1001 0.24851f
C278 voltage_divider_0/m1_3399_17209# avss 0.094199f
C279 level_shifter_0/out_b multiplexer_0/in_1110 0.012179f
C280 avss voltage_divider_0/m1_3935_14185# 0.092648f
C281 multiplexer_0/in_1100 multiplexer_0/in_1101 0.026434f
C282 vin vtrip[1] 0.524944f
C283 avss voltage_divider_0/m1_7155_12295# 0.092648f
C284 vin level_shifter_1/out 0.391713f
C285 multiplexer_0/in_0001 multiplexer_0/in_0100 0.374891f
C286 avss voltage_divider_0/m1_3935_6625# 0.092648f
C287 multiplexer_0/in_1011 avdd 0.18704f
C288 avss voltage_divider_0/m1_3399_577# 0.079556f
C289 avss voltage_divider_0/m1_179_16831# 0.092648f
C290 avss voltage_divider_0/m1_3935_8893# 0.092648f
C291 level_shifter_0/out_b level_shifter_2/out_b 0.128916f
C292 level_shifter_0/out multiplexer_0/trans_gate_m_28/in 0.01094f
C293 avss voltage_divider_0/m1_7155_10783# 0.092648f
C294 avss voltage_divider_0/m1_179_10783# 0.092648f
C295 avss multiplexer_0/trans_gate_m_32/in 0.700225f
C296 level_shifter_1/out multiplexer_0/trans_gate_m_33/in 0.190715f
C297 voltage_divider_0/m1_7691_13807# avss 0.092648f
C298 level_shifter_0/out level_shifter_1/out_b 0.126567f
C299 multiplexer_0/in_1111 multiplexer_0/in_1101 0.471067f
C300 level_shifter_0/out avss 11.112308f
C301 multiplexer_0/in_0101 avss 1.382986f
C302 voltage_divider_0/m1_179_5491# avss 0.092648f
C303 multiplexer_0/trans_gate_m_20/in avdd 0.110125f
C304 voltage_divider_0/m1_7155_16831# avss 0.094199f
C305 vin ena 0.499177f
C306 level_shifter_3/out level_shifter_2/out_b 0.212599f
C307 vin vbg 1.234809f
C308 dvdd vtrip[3] 0.431168f
C309 level_shifter_3/out multiplexer_0/trans_gate_m_34/in 0.851625f
C310 avss multiplexer_0/trans_gate_m_23/in 0.872954f
C311 ibias ena 0.097775f
C312 voltage_divider_0/m1_7691_10027# avss 0.092648f
C313 multiplexer_0/in_0100 multiplexer_0/in_0010 0.018099f
C314 avss voltage_divider_0/m1_179_9271# 0.092648f
C315 level_shifter_0/out multiplexer_0/in_1011 0.072266f
C316 vin avdd 0.915609f
C317 avss voltage_divider_0/m1_3399_3601# 0.079556f
C318 level_shifter_1/in_b vtrip[2] 0.09822f
C319 multiplexer_0/in_0001 avss 1.348022f
C320 avss multiplexer_0/in_1100 0.739738f
C321 initials_0/m4_1419_2382# vin 0.033767f
C322 voltage_divider_0/m1_7155_11539# avss 0.092648f
C323 ibias avdd 0.103351f
C324 avss voltage_divider_0/m1_3399_1333# 0.079556f
C325 multiplexer_0/trans_gate_m_33/in avdd 0.275928f
C326 avss voltage_divider_0/m1_7155_3601# 0.092791f
C327 initials_0/m4_3195_879# initials_0/m4_3195_2379# 0.013296f
C328 avss voltage_divider_0/m1_7155_9271# 0.092648f
C329 voltage_divider_0/m1_10901_199# avss 0.195336f
C330 level_shifter_0/out multiplexer_0/trans_gate_m_20/in 0.039202f
C331 level_shifter_3/out_b level_shifter_2/out 0.167536f
C332 avss multiplexer_0/trans_gate_m_3/out 0.664295f
C333 avss voltage_divider_0/m1_7155_14563# 0.092648f
C334 multiplexer_0/in_1111 avss 0.854435f
C335 voltage_divider_0/m1_7155_17209# avss 0.079556f
C336 multiplexer_0/in_1011 multiplexer_0/in_1100 0.172788f
C337 vin comp_hyst_0/net1 0.334857f
C338 avss voltage_divider_0/m1_3399_4357# 0.092648f
C339 vtrip[2] level_shifter_2/in_b 0.165888f
C340 avss voltage_divider_0/m1_179_8515# 0.092648f
C341 avss multiplexer_0/in_0010 1.622075f
C342 level_shifter_2/out_b multiplexer_0/trans_gate_m_34/in 0.226916f
C343 multiplexer_0/in_0110 multiplexer_0/in_0000 0.01504f
C344 multiplexer_0/trans_gate_m_28/in level_shifter_0/out_b 0.315174f
C345 level_shifter_0/out ibias 0.029237f
C346 vtrip[0] vtrip[3] 0.585874f
C347 level_shifter_0/out multiplexer_0/trans_gate_m_33/in 0.235157f
C348 voltage_divider_0/m1_7155_13051# avss 0.092648f
C349 avss vtrip[3] 1.817329f
C350 avss voltage_divider_0/m1_179_13807# 0.092648f
C351 avss voltage_divider_0/m1_3399_15697# 0.092648f
C352 level_shifter_1/out_b level_shifter_0/out_b 0.148366f
C353 level_shifter_0/out_b avss 9.199488f
C354 multiplexer_0/in_1110 multiplexer_0/in_1101 0.38642f
C355 level_shifter_1/in_b vtrip[1] 0.124413f
C356 avss voltage_divider_0/m1_3399_8137# 0.092648f
C357 multiplexer_0/trans_gate_m_5/out avss 0.719307f
C358 multiplexer_0/in_0000 avdd 0.074544f
C359 voltage_divider_0/m1_7155_6247# avss 0.091766f
C360 level_shifter_3/out level_shifter_1/out_b 0.312288f
C361 level_shifter_3/out avss 3.980763f
C362 voltage_divider_0/m1_179_14563# avss 0.092648f
C363 multiplexer_0/in_1011 level_shifter_0/out_b 0.063584f
C364 vtrip[2] vtrip[1] 2.749246f
C365 level_shifter_1/out level_shifter_2/out 0.127214f
C366 multiplexer_0/in_0110 multiplexer_0/in_0011 1.276962f
C367 level_shifter_3/in_b vtrip[2] 0.161794f
C368 level_shifter_1/in_b ena 0.018249f
C369 voltage_divider_0/m1_7691_16075# avss 0.092648f
C370 level_shifter_2/in_b vtrip[1] 0.151593f
C371 voltage_divider_0/m1_3399_7381# avss 0.092648f
C372 voltage_divider_0/m1_179_4735# avss 0.092648f
C373 multiplexer_0/in_0111 avss 0.927663f
C374 multiplexer_0/in_1110 avss 0.954106f
C375 multiplexer_0/in_1000 multiplexer_0/in_1010 0.488765f
C376 vtrip[2] ena 0.366221f
C377 level_shifter_1/in_b avdd 0.084148f
C378 rocket_0/m1_n9_n9# rocket_0/0 8.528369f
C379 comp_hyst_0/net3 rocket_0/0 20.262209f
C380 comp_hyst_0/net1 rocket_0/0 2.096757f
C381 comp_hyst_0/net4 rocket_0/0 11.427585f
C382 vbg rocket_0/0 11.375807f
C383 ovout rocket_0/0 2.595758f
C384 ibias rocket_0/0 3.449671f
C385 comp_hyst_0/net5 rocket_0/0 31.673025f
C386 comp_hyst_0/ena_b rocket_0/0 9.371887f
C387 dvdd rocket_0/0 0.88126p
C388 ena rocket_0/0 18.616652f
C389 comp_hyst_0/net2 rocket_0/0 7.819766f
C390 initials_0/m4_3195_879# rocket_0/0 0.84996f
C391 initials_0/m4_2307_879# rocket_0/0 0.616607f
C392 initials_0/m4_1419_879# rocket_0/0 0.840328f
C393 initials_0/m4_3395_1229# rocket_0/0 0.590001f
C394 initials_0/m4_2374_1229# rocket_0/0 0.58922f
C395 initials_0/m4_1419_1229# rocket_0/0 0.668524f
C396 initials_0/m4_3195_2379# rocket_0/0 1.075676f
C397 initials_0/m4_2474_2379# rocket_0/0 0.533313f
C398 initials_0/m4_1419_2382# rocket_0/0 1.186582f
C399 vtrip[3] rocket_0/0 5.541124f
C400 level_shifter_3/in_b rocket_0/0 3.086004f
C401 vtrip[2] rocket_0/0 5.494162f
C402 level_shifter_2/in_b rocket_0/0 3.059048f
C403 vtrip[1] rocket_0/0 5.858896f
C404 level_shifter_1/in_b rocket_0/0 3.082257f
C405 vtrip[0] rocket_0/0 6.905421f
C406 level_shifter_0/in_b rocket_0/0 3.041645f
C407 level_shifter_1/out rocket_0/0 10.188188f
C408 multiplexer_0/in_1100 rocket_0/0 2.538941f
C409 multiplexer_0/trans_gate_m_20/in rocket_0/0 1.350471f
C410 level_shifter_1/out_b rocket_0/0 8.553854f
C411 multiplexer_0/trans_gate_m_37/in rocket_0/0 1.382917f
C412 level_shifter_0/out rocket_0/0 18.046806f
C413 multiplexer_0/trans_gate_m_9/out rocket_0/0 1.746898f
C414 multiplexer_0/in_1101 rocket_0/0 2.635137f
C415 level_shifter_0/out_b rocket_0/0 17.55795f
C416 multiplexer_0/trans_gate_m_33/in rocket_0/0 1.978841f
C417 multiplexer_0/in_1111 rocket_0/0 3.21071f
C418 level_shifter_2/out rocket_0/0 3.723293f
C419 multiplexer_0/trans_gate_m_34/in rocket_0/0 1.978869f
C420 level_shifter_2/out_b rocket_0/0 4.578737f
C421 avdd rocket_0/0 0.901897p
C422 multiplexer_0/in_0000 rocket_0/0 3.032357f
C423 multiplexer_0/trans_gate_m_7/out rocket_0/0 1.144867f
C424 multiplexer_0/in_1110 rocket_0/0 3.046156f
C425 multiplexer_0/trans_gate_m_28/in rocket_0/0 1.129369f
C426 multiplexer_0/trans_gate_m_31/in rocket_0/0 1.774978f
C427 multiplexer_0/in_0001 rocket_0/0 2.865136f
C428 multiplexer_0/in_1010 rocket_0/0 2.823186f
C429 multiplexer_0/in_0100 rocket_0/0 3.018654f
C430 multiplexer_0/trans_gate_m_5/out rocket_0/0 1.147648f
C431 multiplexer_0/in_1011 rocket_0/0 2.58388f
C432 level_shifter_3/out rocket_0/0 3.05246f
C433 vin rocket_0/0 17.129452f
C434 level_shifter_3/out_b rocket_0/0 3.434802f
C435 multiplexer_0/trans_gate_m_27/in rocket_0/0 1.810418f
C436 multiplexer_0/in_0101 rocket_0/0 2.888583f
C437 multiplexer_0/trans_gate_m_3/out rocket_0/0 1.147648f
C438 multiplexer_0/in_0111 rocket_0/0 2.841224f
C439 multiplexer_0/trans_gate_m_23/in rocket_0/0 1.808818f
C440 multiplexer_0/in_1001 rocket_0/0 2.53703f
C441 multiplexer_0/in_0110 rocket_0/0 2.925628f
C442 multiplexer_0/trans_gate_m_32/in rocket_0/0 1.133956f
C443 multiplexer_0/in_1000 rocket_0/0 2.728564f
C444 multiplexer_0/trans_gate_m_29/in rocket_0/0 1.137561f
C445 multiplexer_0/in_0011 rocket_0/0 2.839224f
C446 multiplexer_0/in_0010 rocket_0/0 3.499047f
C447 voltage_divider_0/m1_10911_16453# rocket_0/0 0.789952f
C448 voltage_divider_0/m1_7691_16075# rocket_0/0 0.600369f
C449 voltage_divider_0/m1_10911_15697# rocket_0/0 0.789096f
C450 voltage_divider_0/m1_7691_15319# rocket_0/0 0.599493f
C451 voltage_divider_0/m1_10911_14941# rocket_0/0 0.789055f
C452 voltage_divider_0/m1_7691_14563# rocket_0/0 0.599493f
C453 voltage_divider_0/m1_10911_14185# rocket_0/0 0.789055f
C454 voltage_divider_0/m1_7691_13807# rocket_0/0 0.599493f
C455 voltage_divider_0/m1_10911_13429# rocket_0/0 0.789055f
C456 voltage_divider_0/m1_7691_13051# rocket_0/0 0.599493f
C457 voltage_divider_0/m1_10911_12673# rocket_0/0 0.789055f
C458 voltage_divider_0/m1_7691_12295# rocket_0/0 0.599493f
C459 voltage_divider_0/m1_10911_11917# rocket_0/0 0.789055f
C460 voltage_divider_0/51 rocket_0/0 0.599493f
C461 voltage_divider_0/m1_7691_10783# rocket_0/0 0.599493f
C462 voltage_divider_0/m1_7691_10027# rocket_0/0 0.599493f
C463 voltage_divider_0/m1_7691_9271# rocket_0/0 0.599493f
C464 voltage_divider_0/m1_10901_8137# rocket_0/0 0.800173f
C465 voltage_divider_0/m1_7691_7003# rocket_0/0 0.599493f
C466 voltage_divider_0/m1_10911_2845# rocket_0/0 0.789055f
C467 voltage_divider_0/m1_10911_2089# rocket_0/0 0.789055f
C468 voltage_divider_0/m1_10911_1333# rocket_0/0 0.789096f
C469 voltage_divider_0/m1_10911_577# rocket_0/0 0.791315f
C470 voltage_divider_0/m1_10901_199# rocket_0/0 3.463708f
C471 voltage_divider_0/m1_7155_17209# rocket_0/0 0.883249f
C472 voltage_divider_0/m1_7155_16831# rocket_0/0 0.604193f
C473 voltage_divider_0/m1_3935_16453# rocket_0/0 0.601754f
C474 voltage_divider_0/m1_7155_16075# rocket_0/0 0.600369f
C475 voltage_divider_0/m1_3935_15697# rocket_0/0 0.599535f
C476 voltage_divider_0/m1_7155_15319# rocket_0/0 0.599493f
C477 voltage_divider_0/m1_3935_14941# rocket_0/0 0.599493f
C478 voltage_divider_0/m1_7155_14563# rocket_0/0 0.599493f
C479 voltage_divider_0/m1_3935_14185# rocket_0/0 0.599493f
C480 voltage_divider_0/m1_7155_13807# rocket_0/0 0.599493f
C481 voltage_divider_0/m1_3935_13429# rocket_0/0 0.599493f
C482 voltage_divider_0/m1_7155_13051# rocket_0/0 0.599493f
C483 voltage_divider_0/m1_3935_12673# rocket_0/0 0.599493f
C484 voltage_divider_0/m1_7155_12295# rocket_0/0 0.599493f
C485 voltage_divider_0/m1_3935_11917# rocket_0/0 0.599493f
C486 voltage_divider_0/m1_7155_11539# rocket_0/0 0.599493f
C487 voltage_divider_0/m1_3935_11161# rocket_0/0 0.599493f
C488 voltage_divider_0/m1_7155_10783# rocket_0/0 0.599493f
C489 voltage_divider_0/m1_3935_10405# rocket_0/0 0.599493f
C490 voltage_divider_0/m1_7155_10027# rocket_0/0 0.599493f
C491 voltage_divider_0/m1_3935_9649# rocket_0/0 0.599493f
C492 voltage_divider_0/m1_7155_9271# rocket_0/0 0.599493f
C493 voltage_divider_0/m1_3935_8893# rocket_0/0 0.599493f
C494 voltage_divider_0/m1_7155_8515# rocket_0/0 0.598612f
C495 voltage_divider_0/m1_3935_8137# rocket_0/0 0.599493f
C496 voltage_divider_0/m1_7155_7759# rocket_0/0 0.598612f
C497 voltage_divider_0/m1_3935_7381# rocket_0/0 0.599493f
C498 voltage_divider_0/m1_7155_7003# rocket_0/0 0.599493f
C499 voltage_divider_0/m1_3935_6625# rocket_0/0 0.599493f
C500 voltage_divider_0/m1_7155_6247# rocket_0/0 0.598612f
C501 voltage_divider_0/m1_3935_5869# rocket_0/0 0.599493f
C502 voltage_divider_0/m1_7155_5491# rocket_0/0 0.598612f
C503 voltage_divider_0/m1_3935_5113# rocket_0/0 0.599493f
C504 voltage_divider_0/m1_7155_4735# rocket_0/0 0.598612f
C505 voltage_divider_0/m1_3935_4357# rocket_0/0 0.599493f
C506 voltage_divider_0/m1_7155_3979# rocket_0/0 0.598612f
C507 voltage_divider_0/m1_7155_3601# rocket_0/0 0.599576f
C508 voltage_divider_0/m1_7155_3223# rocket_0/0 0.583453f
C509 voltage_divider_0/m1_7155_2845# rocket_0/0 0.583453f
C510 voltage_divider_0/m1_7155_2467# rocket_0/0 0.583453f
C511 voltage_divider_0/m1_7155_2089# rocket_0/0 0.583453f
C512 voltage_divider_0/m1_7155_1711# rocket_0/0 0.583453f
C513 voltage_divider_0/m1_7155_1333# rocket_0/0 0.583545f
C514 voltage_divider_0/m1_7155_955# rocket_0/0 0.584937f
C515 voltage_divider_0/m1_7155_577# rocket_0/0 0.586355f
C516 voltage_divider_0/m1_7155_199# rocket_0/0 0.883249f
C517 voltage_divider_0/m1_3399_17209# rocket_0/0 0.901087f
C518 voltage_divider_0/m1_179_16831# rocket_0/0 0.924812f
C519 voltage_divider_0/m1_3399_16453# rocket_0/0 0.601754f
C520 voltage_divider_0/m1_179_16075# rocket_0/0 0.78993f
C521 voltage_divider_0/m1_3399_15697# rocket_0/0 0.599535f
C522 voltage_divider_0/m1_179_15319# rocket_0/0 0.789055f
C523 voltage_divider_0/m1_3399_14941# rocket_0/0 0.599493f
C524 voltage_divider_0/m1_179_14563# rocket_0/0 0.789055f
C525 voltage_divider_0/m1_3399_14185# rocket_0/0 0.599493f
C526 voltage_divider_0/m1_179_13807# rocket_0/0 0.789055f
C527 voltage_divider_0/m1_3399_13429# rocket_0/0 0.599493f
C528 voltage_divider_0/m1_179_13051# rocket_0/0 0.789055f
C529 voltage_divider_0/m1_3399_12673# rocket_0/0 0.599493f
C530 voltage_divider_0/m1_179_12295# rocket_0/0 0.789055f
C531 voltage_divider_0/m1_3399_11917# rocket_0/0 0.599493f
C532 voltage_divider_0/m1_179_11539# rocket_0/0 0.789055f
C533 voltage_divider_0/m1_3399_11161# rocket_0/0 0.599493f
C534 voltage_divider_0/m1_179_10783# rocket_0/0 0.789055f
C535 voltage_divider_0/m1_3399_10405# rocket_0/0 0.599493f
C536 voltage_divider_0/m1_179_10027# rocket_0/0 0.789055f
C537 voltage_divider_0/m1_3399_9649# rocket_0/0 0.599493f
C538 voltage_divider_0/m1_179_9271# rocket_0/0 0.789055f
C539 voltage_divider_0/m1_3399_8893# rocket_0/0 0.599493f
C540 voltage_divider_0/m1_179_8515# rocket_0/0 0.789055f
C541 voltage_divider_0/m1_3399_8137# rocket_0/0 0.599493f
C542 voltage_divider_0/m1_179_7759# rocket_0/0 0.789055f
C543 voltage_divider_0/m1_3399_7381# rocket_0/0 0.599493f
C544 voltage_divider_0/m1_179_7003# rocket_0/0 0.789055f
C545 voltage_divider_0/m1_3399_6625# rocket_0/0 0.599493f
C546 voltage_divider_0/m1_179_6247# rocket_0/0 0.789055f
C547 voltage_divider_0/m1_3399_5869# rocket_0/0 0.599493f
C548 voltage_divider_0/m1_179_5491# rocket_0/0 0.789055f
C549 voltage_divider_0/m1_3399_5113# rocket_0/0 0.599493f
C550 voltage_divider_0/m1_179_4735# rocket_0/0 0.789055f
C551 voltage_divider_0/m1_3399_4357# rocket_0/0 0.599493f
C552 voltage_divider_0/m1_3399_3979# rocket_0/0 0.601291f
C553 voltage_divider_0/m1_179_3979# rocket_0/0 0.789055f
C554 voltage_divider_0/m1_3399_3601# rocket_0/0 0.583453f
C555 voltage_divider_0/m1_3399_3223# rocket_0/0 0.583453f
C556 voltage_divider_0/m1_179_3223# rocket_0/0 0.789055f
C557 voltage_divider_0/m1_3399_2845# rocket_0/0 0.583453f
C558 voltage_divider_0/m1_3399_2467# rocket_0/0 0.583453f
C559 voltage_divider_0/m1_179_2467# rocket_0/0 0.789055f
C560 voltage_divider_0/m1_3399_2089# rocket_0/0 0.583453f
C561 voltage_divider_0/m1_3399_1711# rocket_0/0 0.583453f
C562 voltage_divider_0/m1_179_1711# rocket_0/0 0.789055f
C563 voltage_divider_0/m1_3399_1333# rocket_0/0 0.583545f
C564 voltage_divider_0/m1_3399_955# rocket_0/0 0.584937f
C565 voltage_divider_0/m1_179_955# rocket_0/0 0.78993f
C566 voltage_divider_0/m1_3399_577# rocket_0/0 0.586355f
C567 voltage_divider_0/m1_3399_199# rocket_0/0 0.883249f
C568 voltage_divider_0/m1_179_199# rocket_0/0 0.924812f
.ends


magic
tech sky130A
magscale 1 2
timestamp 1712948219
<< nwell >>
rect 15899 1815 15954 1823
rect 14281 1580 15936 1584
rect 14281 1577 15921 1580
rect 15918 1505 15921 1577
<< pwell >>
rect 14055 -5363 14471 -4997
<< locali >>
rect 1703 2440 13650 2528
rect 1703 2216 1864 2440
rect 13550 2216 13650 2440
rect 1703 1464 13650 2216
rect 13167 -698 13650 1464
rect 6914 -1024 13167 -698
rect 8720 -1590 9046 -1024
rect 9966 -1590 10292 -1024
rect 12212 -1590 12648 -1024
rect 6914 -1915 8568 -1590
rect 6914 -2007 7208 -1915
rect 9968 -2294 10292 -1786
rect 9048 -2334 10292 -2294
rect 12212 -2334 12648 -2134
rect 9048 -2512 12648 -2334
rect 9048 -3060 9398 -2512
rect 12090 -3060 12648 -2512
rect 9048 -3082 12648 -3060
rect 13168 -3082 13663 -2133
rect 9048 -3298 13663 -3082
rect 6845 -4109 7205 -3821
rect 7139 -4453 7205 -4109
rect 6845 -4533 7205 -4453
rect 8565 -4360 9048 -3820
rect 13368 -4360 13663 -3298
rect 8565 -4533 13663 -4360
rect 6845 -4967 13663 -4533
rect 6845 -5028 16899 -4967
rect 6845 -5252 6970 -5028
rect 13292 -5033 16899 -5028
rect 13292 -5252 14091 -5033
rect 6845 -5327 14091 -5252
rect 14435 -5327 16128 -5033
rect 16472 -5327 16899 -5033
<< viali >>
rect 1864 2216 13550 2440
rect 6970 -5252 13292 -5028
<< metal1 >>
rect 1703 2440 13650 2528
rect 1703 2216 1864 2440
rect 13550 2432 13650 2440
rect 13550 2386 16434 2432
rect 13550 2216 13650 2386
rect 1703 2135 13650 2216
rect 1702 1804 13650 2135
rect 1702 1796 13404 1804
rect 1702 1608 2205 1796
rect 2425 1608 5688 1796
rect 5908 1608 9176 1796
rect 9396 1616 13404 1796
rect 13624 1616 13650 1804
rect 9396 1608 13650 1616
rect 1702 1544 13650 1608
rect 13758 2104 13804 2386
rect 14016 2104 14062 2386
rect 14190 2104 14290 2386
rect 15902 2104 15948 2386
rect 16130 2104 16176 2386
rect 16388 2104 16434 2386
rect 13758 2058 16434 2104
rect 13758 1900 13804 2058
rect 14016 1900 14062 2058
rect 13758 1854 13822 1900
rect 14001 1854 14062 1900
rect 14286 1861 14296 1918
rect 15896 1861 15906 1918
rect 14286 1854 15906 1861
rect 16130 1900 16176 2058
rect 16388 1900 16434 2058
rect 16130 1854 16199 1900
rect 16374 1854 16434 1900
rect 13758 1572 13804 1854
rect 14016 1572 14062 1854
rect 1811 1368 1857 1544
rect 5555 1368 5829 1544
rect 9041 1368 9315 1544
rect 13013 1368 13059 1544
rect 1811 1322 13059 1368
rect 1811 1040 1857 1322
rect 2069 1040 2115 1322
rect 2265 1040 2343 1322
rect 5555 1040 5601 1322
rect 5751 1040 5829 1322
rect 9041 1040 9087 1322
rect 9237 1040 9315 1322
rect 12527 1040 12573 1322
rect 12755 1040 12801 1322
rect 13013 1040 13059 1322
rect 1811 994 13059 1040
rect 1811 836 1857 994
rect 2069 836 2115 994
rect 1811 790 1888 836
rect 2051 790 2115 836
rect 2339 797 2349 853
rect 5549 797 5559 853
rect 2339 790 5559 797
rect 5825 797 5835 853
rect 9035 797 9087 853
rect 5825 790 9087 797
rect 9311 797 9321 853
rect 12521 797 12531 853
rect 9311 790 12531 797
rect 12755 836 12801 994
rect 13013 836 13059 994
rect 12755 790 12830 836
rect 12992 790 13059 836
rect 1811 508 1857 790
rect 2069 508 2115 790
rect 9041 749 9087 790
rect 1811 462 1884 508
rect 2053 462 2115 508
rect 1811 304 1857 462
rect 2069 304 2115 462
rect 1811 258 1885 304
rect 2056 258 2115 304
rect 1811 -24 1857 258
rect 2069 -24 2115 258
rect 2265 549 2291 749
rect 2343 549 2353 749
rect 5545 549 5555 749
rect 5607 549 5617 749
rect 5751 549 5777 749
rect 5829 549 5839 749
rect 9237 549 9263 749
rect 9315 549 9325 749
rect 12517 549 12527 749
rect 12579 549 12589 749
rect 2265 17 2311 549
rect 2339 501 5559 508
rect 2339 445 2349 501
rect 5549 445 5559 501
rect 2339 265 2349 321
rect 5549 265 5559 321
rect 2339 258 5559 265
rect 5545 17 5555 217
rect 5607 17 5617 217
rect 5751 17 5797 549
rect 9041 508 9087 549
rect 5825 501 9087 508
rect 5825 445 5835 501
rect 9035 445 9087 501
rect 5825 265 5835 321
rect 9035 265 9087 321
rect 5825 258 9087 265
rect 9041 217 9087 258
rect 9237 17 9283 549
rect 12755 508 12801 790
rect 13013 508 13059 790
rect 13758 1526 13826 1572
rect 14004 1526 14062 1572
rect 13758 1368 13804 1526
rect 14016 1368 14062 1526
rect 13758 1322 13826 1368
rect 14004 1322 14062 1368
rect 13758 1040 13804 1322
rect 14016 1040 14062 1322
rect 13758 994 13828 1040
rect 14004 994 14062 1040
rect 13758 836 13804 994
rect 14016 836 14062 994
rect 13758 790 13824 836
rect 13994 790 14062 836
rect 13758 508 13804 790
rect 14016 508 14062 790
rect 9311 501 12531 508
rect 9311 445 9321 501
rect 12521 445 12531 501
rect 12755 462 12831 508
rect 12995 462 13826 508
rect 14003 462 14062 508
rect 9311 265 9321 321
rect 12521 265 12531 321
rect 9311 258 12531 265
rect 12755 304 12801 462
rect 13013 304 13804 462
rect 14016 304 14062 462
rect 12755 258 12829 304
rect 12993 258 13822 304
rect 14001 258 14062 304
rect 12517 17 12527 217
rect 12579 17 12589 217
rect 9041 -24 9087 17
rect 12755 -24 12801 258
rect 13013 -24 13059 258
rect 1811 -70 1889 -24
rect 2052 -70 2115 -24
rect 1811 -228 1857 -70
rect 2069 -228 2115 -70
rect 2339 -31 5559 -24
rect 2339 -87 2349 -31
rect 5549 -87 5559 -31
rect 5825 -31 9087 -24
rect 5825 -87 5835 -31
rect 9035 -87 9087 -31
rect 9311 -31 12531 -24
rect 9311 -87 9321 -31
rect 12521 -87 12531 -31
rect 12755 -70 12834 -24
rect 12990 -70 13059 -24
rect 12755 -228 12801 -70
rect 13013 -228 13059 -70
rect 1811 -274 13059 -228
rect 1811 -556 1857 -274
rect 2069 -556 2115 -274
rect 2265 -556 2343 -274
rect 5555 -556 5601 -274
rect 5751 -556 5829 -274
rect 9041 -556 9087 -274
rect 9237 -556 9315 -274
rect 12527 -556 12573 -274
rect 12755 -556 12801 -274
rect 13013 -556 13059 -274
rect 13758 -24 13804 258
rect 14016 -24 14062 258
rect 14190 1613 14238 1813
rect 14290 1613 14300 1813
rect 15892 1613 15902 1813
rect 15954 1613 15964 1813
rect 14190 17 14258 1613
rect 16130 1572 16176 1854
rect 16388 1572 16434 1854
rect 14286 1565 15906 1572
rect 14286 1508 14296 1565
rect 15896 1508 15906 1565
rect 16130 1526 16200 1572
rect 16377 1526 16434 1572
rect 14286 1329 14296 1386
rect 15896 1329 15948 1386
rect 14286 1322 15948 1329
rect 15902 1280 15948 1322
rect 16130 1368 16176 1526
rect 16388 1368 16434 1526
rect 16130 1322 16194 1368
rect 16375 1322 16434 1368
rect 15902 1040 15948 1081
rect 14287 1033 15948 1040
rect 14287 976 14297 1033
rect 15897 976 15948 1033
rect 16130 1040 16176 1322
rect 16388 1040 16434 1322
rect 16130 994 16197 1040
rect 16375 994 16434 1040
rect 14286 797 14296 854
rect 15896 797 15948 854
rect 14286 790 15948 797
rect 15902 749 15948 790
rect 16130 836 16176 994
rect 16388 836 16434 994
rect 16130 790 16198 836
rect 16374 790 16434 836
rect 15902 508 15948 549
rect 14286 501 15948 508
rect 14286 444 14296 501
rect 15896 444 15948 501
rect 16130 508 16176 790
rect 16388 508 16434 790
rect 16130 462 16198 508
rect 16376 462 16434 508
rect 14286 265 14296 322
rect 15896 265 15906 322
rect 14286 258 15906 265
rect 16130 304 16176 462
rect 16388 304 16434 462
rect 16130 258 16195 304
rect 16370 258 16434 304
rect 15892 17 15902 217
rect 15954 17 15964 217
rect 16130 -24 16176 258
rect 16388 -24 16434 258
rect 13758 -70 13824 -24
rect 13998 -70 14062 -24
rect 13758 -228 13804 -70
rect 14016 -228 14062 -70
rect 14286 -31 15906 -24
rect 14286 -88 14296 -31
rect 15896 -88 15906 -31
rect 16130 -70 16200 -24
rect 16367 -70 16434 -24
rect 16130 -228 16176 -70
rect 16388 -228 16434 -70
rect 13758 -274 16434 -228
rect 13758 -556 13804 -274
rect 14016 -556 14062 -274
rect 14190 -556 14291 -274
rect 15902 -556 15948 -274
rect 16130 -556 16176 -274
rect 16388 -556 16434 -274
rect 1811 -602 16434 -556
rect 6948 -1207 7036 -602
rect 7064 -1159 7074 -1107
rect 7674 -1159 7684 -1107
rect 7834 -1207 7922 -602
rect 7950 -1159 7960 -1107
rect 8560 -1159 8570 -1107
rect 9080 -1207 9168 -602
rect 9196 -1159 9206 -1107
rect 9806 -1159 9816 -1107
rect 10326 -1207 10414 -602
rect 10442 -1159 10452 -1107
rect 12052 -1159 12062 -1107
rect 12682 -1207 12770 -602
rect 13328 -1017 16661 -839
rect 12798 -1159 12808 -1107
rect 13008 -1159 13018 -1107
rect 13328 -1206 13505 -1017
rect 13092 -1207 13505 -1206
rect 6948 -1407 7068 -1207
rect 7670 -1407 7680 -1207
rect 7732 -1407 7742 -1207
rect 6948 -1915 7036 -1407
rect 7834 -1411 7948 -1207
rect 8556 -1407 8566 -1207
rect 8618 -1407 8628 -1207
rect 9080 -1407 9200 -1207
rect 9812 -1407 9890 -1207
rect 10326 -1407 10446 -1207
rect 12048 -1407 12058 -1207
rect 12110 -1407 12120 -1207
rect 7064 -1507 7074 -1455
rect 7674 -1507 7684 -1455
rect 7950 -1507 7960 -1455
rect 8560 -1507 8570 -1455
rect 9196 -1507 9206 -1455
rect 9806 -1507 9816 -1455
rect 9844 -1643 9890 -1407
rect 10442 -1507 10452 -1455
rect 12052 -1507 12062 -1455
rect 9128 -1689 9890 -1643
rect 6948 -2007 7292 -1915
rect 9128 -1920 9174 -1689
rect 12682 -1807 12802 -1207
rect 13014 -1383 13505 -1207
rect 16725 -1309 16771 -1308
rect 13791 -1355 16771 -1309
rect 13014 -1384 13504 -1383
rect 13014 -1807 13134 -1384
rect 9202 -1872 9212 -1820
rect 9808 -1872 9818 -1820
rect 10400 -1912 10452 -1860
rect 12052 -1912 12062 -1860
rect 12798 -1907 12808 -1855
rect 13008 -1907 13018 -1855
rect 9128 -2120 9150 -1920
rect 9202 -2120 9212 -1920
rect 9814 -2120 9934 -1920
rect 10400 -1928 10480 -1912
rect 10400 -1960 10446 -1928
rect 9198 -2220 9208 -2168
rect 9804 -2220 9814 -2168
rect 9842 -2372 9934 -2120
rect 10384 -2160 10394 -1960
rect 10446 -2160 10456 -1960
rect 12060 -2160 12178 -1960
rect 13046 -2026 13134 -1807
rect 10400 -2192 10446 -2160
rect 10400 -2208 10478 -2192
rect 10400 -2260 10452 -2208
rect 12052 -2260 12062 -2208
rect 12090 -2372 12178 -2160
rect 9842 -2464 12178 -2372
rect 12682 -2098 13134 -2026
rect 13791 -1619 13837 -1355
rect 14049 -1619 14095 -1355
rect 14429 -1619 14475 -1355
rect 16087 -1619 16133 -1355
rect 16467 -1619 16513 -1355
rect 16725 -1619 16771 -1355
rect 13791 -1665 16771 -1619
rect 13791 -1895 13837 -1665
rect 14049 -1895 14095 -1665
rect 13791 -1941 13854 -1895
rect 14038 -1941 14095 -1895
rect 14471 -1925 14481 -1873
rect 16081 -1925 16091 -1873
rect 14471 -1941 16091 -1925
rect 16467 -1895 16513 -1665
rect 16725 -1895 16771 -1665
rect 16467 -1941 16530 -1895
rect 16710 -1941 16771 -1895
rect 12682 -2308 12770 -2098
rect 12798 -2260 12808 -2208
rect 13008 -2260 13018 -2208
rect 13791 -2265 13837 -1941
rect 14049 -2265 14095 -1941
rect 14413 -2233 14423 -1973
rect 14475 -2233 14485 -1973
rect 9556 -2638 9566 -2586
rect 10166 -2638 10176 -2586
rect 10204 -2686 10284 -2464
rect 10442 -2638 10452 -2586
rect 11052 -2638 11062 -2586
rect 11090 -2686 11170 -2464
rect 11328 -2638 11338 -2586
rect 11938 -2638 11948 -2586
rect 11976 -2686 12056 -2464
rect 9498 -2886 9508 -2686
rect 9560 -2886 9570 -2686
rect 10164 -2886 10284 -2686
rect 10384 -2886 10394 -2686
rect 10446 -2886 10456 -2686
rect 11050 -2886 11170 -2686
rect 11270 -2886 11280 -2686
rect 11332 -2886 11342 -2686
rect 11936 -2886 12056 -2686
rect 9556 -2986 9566 -2934
rect 10166 -2986 10176 -2934
rect 10204 -3129 10284 -2886
rect 10442 -2986 10452 -2934
rect 11052 -2986 11062 -2934
rect 11090 -3126 11170 -2886
rect 11328 -2986 11338 -2934
rect 11938 -2986 11948 -2934
rect 11976 -3126 12056 -2886
rect 12682 -2908 12750 -2308
rect 12802 -2908 12812 -2308
rect 13014 -2908 13134 -2308
rect 12798 -3008 12808 -2956
rect 13008 -3008 13018 -2956
rect 13046 -3126 13134 -2908
rect 13791 -2311 13853 -2265
rect 14031 -2311 14095 -2265
rect 13791 -2541 13837 -2311
rect 14049 -2541 14095 -2311
rect 14471 -2281 16091 -2265
rect 14471 -2333 14481 -2281
rect 16081 -2333 16091 -2281
rect 13791 -2587 13854 -2541
rect 14032 -2587 14095 -2541
rect 14471 -2571 14481 -2519
rect 16081 -2571 16091 -2519
rect 14471 -2587 16091 -2571
rect 13791 -2911 13837 -2587
rect 14049 -2911 14095 -2587
rect 14413 -2879 14423 -2619
rect 14475 -2879 14485 -2619
rect 13791 -2957 13847 -2911
rect 14038 -2957 14095 -2911
rect 13791 -3126 13837 -2957
rect 11090 -3129 13837 -3126
rect 10204 -3187 13837 -3129
rect 14049 -3187 14095 -2957
rect 14471 -2979 14481 -2927
rect 16081 -2979 16091 -2927
rect 10204 -3206 13850 -3187
rect 10204 -3209 11187 -3206
rect 9140 -3424 9208 -3372
rect 13208 -3424 13218 -3372
rect 9140 -3440 13218 -3424
rect 9140 -3472 9212 -3440
rect 9140 -3672 9150 -3472
rect 9202 -3672 9212 -3472
rect 9140 -3704 9212 -3672
rect 7108 -3786 7206 -3710
rect 9140 -3720 13218 -3704
rect 9140 -3772 9208 -3720
rect 13208 -3772 13218 -3720
rect 9198 -3938 9208 -3886
rect 13208 -3938 13218 -3886
rect 9198 -3954 13218 -3938
rect 9140 -4186 9150 -3986
rect 9202 -4186 9212 -3986
rect 6943 -4351 6953 -4211
rect 7031 -4351 7041 -4211
rect 9198 -4234 13218 -4218
rect 9198 -4286 9208 -4234
rect 13208 -4286 13218 -4234
rect 13246 -4441 13334 -3206
rect 8565 -4479 13334 -4441
rect 13791 -3233 13850 -3206
rect 14037 -3233 14095 -3187
rect 14471 -3217 14481 -3165
rect 16081 -3217 16091 -3165
rect 13791 -3557 13837 -3233
rect 14049 -3557 14095 -3233
rect 14413 -3525 14423 -3265
rect 14475 -3525 14485 -3265
rect 13791 -3603 13852 -3557
rect 14034 -3603 14095 -3557
rect 13791 -3833 13837 -3603
rect 14049 -3833 14095 -3603
rect 14471 -3573 16091 -3557
rect 14471 -3625 14481 -3573
rect 16081 -3625 16091 -3573
rect 13791 -3879 13847 -3833
rect 14038 -3879 14095 -3833
rect 14471 -3863 14481 -3811
rect 16081 -3863 16091 -3811
rect 14471 -3879 16091 -3863
rect 13791 -4203 13837 -3879
rect 14049 -4203 14095 -3879
rect 14413 -4171 14423 -3911
rect 14475 -4171 14485 -3911
rect 13791 -4249 13850 -4203
rect 14037 -4249 14095 -4203
rect 13791 -4479 13837 -4249
rect 14049 -4479 14095 -4249
rect 14471 -4219 16091 -4203
rect 14471 -4271 14481 -4219
rect 16081 -4271 16091 -4219
rect 16119 -4337 16165 -1973
rect 16467 -2265 16513 -1941
rect 16725 -2265 16771 -1941
rect 16467 -2311 16530 -2265
rect 16710 -2311 16771 -2265
rect 16467 -2541 16513 -2311
rect 16725 -2541 16771 -2311
rect 16467 -2587 16529 -2541
rect 16708 -2587 16771 -2541
rect 16467 -2911 16513 -2587
rect 16725 -2911 16771 -2587
rect 16467 -2957 16529 -2911
rect 16712 -2957 16771 -2911
rect 16467 -3187 16513 -2957
rect 16725 -3187 16771 -2957
rect 16467 -3233 16528 -3187
rect 16714 -3233 16771 -3187
rect 16467 -3557 16513 -3233
rect 16725 -3557 16771 -3233
rect 16467 -3603 16527 -3557
rect 16712 -3603 16771 -3557
rect 16467 -3833 16513 -3603
rect 16725 -3833 16771 -3603
rect 16467 -3879 16530 -3833
rect 16710 -3879 16771 -3833
rect 16467 -4203 16513 -3879
rect 16725 -4203 16771 -3879
rect 16467 -4249 16528 -4203
rect 16715 -4249 16771 -4203
rect 16056 -4389 16066 -4337
rect 16206 -4389 16216 -4337
rect 16467 -4479 16513 -4249
rect 16725 -4479 16771 -4249
rect 8565 -4525 16771 -4479
rect 8565 -4533 13837 -4525
rect 6845 -4789 13837 -4533
rect 14049 -4789 14095 -4525
rect 14429 -4789 14475 -4525
rect 16087 -4789 16133 -4525
rect 16467 -4789 16513 -4525
rect 16725 -4789 16771 -4525
rect 6845 -4835 16771 -4789
rect 6845 -5028 13404 -4835
rect 16467 -4836 16513 -4835
rect 6845 -5252 6970 -5028
rect 13292 -5252 13404 -5028
rect 14183 -5219 14193 -5141
rect 14333 -5219 14343 -5141
rect 16221 -5220 16231 -5141
rect 16370 -5220 16380 -5141
rect 6845 -5327 13404 -5252
<< via1 >>
rect 2205 1608 2425 1796
rect 5688 1608 5908 1796
rect 9176 1608 9396 1796
rect 13404 1616 13624 1804
rect 14296 1861 15896 1918
rect 2349 797 5549 853
rect 5835 797 9035 853
rect 9321 797 12521 853
rect 2291 549 2343 749
rect 5555 549 5607 749
rect 5777 549 5829 749
rect 9263 549 9315 749
rect 12527 549 12579 749
rect 2349 445 5549 501
rect 2349 265 5549 321
rect 5555 17 5607 217
rect 5835 445 9035 501
rect 5835 265 9035 321
rect 9321 445 12521 501
rect 9321 265 12521 321
rect 12527 17 12579 217
rect 2349 -87 5549 -31
rect 5835 -87 9035 -31
rect 9321 -87 12521 -31
rect 14238 1613 14290 1813
rect 15902 1613 15954 1813
rect 14296 1508 15896 1565
rect 14296 1329 15896 1386
rect 14297 976 15897 1033
rect 14296 797 15896 854
rect 14296 444 15896 501
rect 14296 265 15896 322
rect 15902 17 15954 217
rect 14296 -88 15896 -31
rect 7074 -1159 7674 -1107
rect 7960 -1159 8560 -1107
rect 9206 -1159 9806 -1107
rect 10452 -1159 12052 -1107
rect 12808 -1159 13008 -1107
rect 7680 -1407 7732 -1207
rect 8566 -1407 8618 -1207
rect 12058 -1407 12110 -1207
rect 7074 -1507 7674 -1455
rect 7960 -1507 8560 -1455
rect 9206 -1507 9806 -1455
rect 10452 -1507 12052 -1455
rect 9212 -1872 9808 -1820
rect 10452 -1912 12052 -1860
rect 12808 -1907 13008 -1855
rect 9150 -2120 9202 -1920
rect 9208 -2220 9804 -2168
rect 10394 -2160 10446 -1960
rect 10452 -2260 12052 -2208
rect 14481 -1925 16081 -1873
rect 12808 -2260 13008 -2208
rect 14423 -2233 14475 -1973
rect 9566 -2638 10166 -2586
rect 10452 -2638 11052 -2586
rect 11338 -2638 11938 -2586
rect 9508 -2886 9560 -2686
rect 10394 -2886 10446 -2686
rect 11280 -2886 11332 -2686
rect 9566 -2986 10166 -2934
rect 10452 -2986 11052 -2934
rect 11338 -2986 11938 -2934
rect 12750 -2908 12802 -2308
rect 12808 -3008 13008 -2956
rect 14481 -2333 16081 -2281
rect 14481 -2571 16081 -2519
rect 14423 -2879 14475 -2619
rect 14481 -2979 16081 -2927
rect 9208 -3424 13208 -3372
rect 9150 -3672 9202 -3472
rect 9208 -3772 13208 -3720
rect 9208 -3938 13208 -3886
rect 9150 -4186 9202 -3986
rect 6953 -4351 7031 -4211
rect 9208 -4286 13208 -4234
rect 14481 -3217 16081 -3165
rect 14423 -3525 14475 -3265
rect 14481 -3625 16081 -3573
rect 14481 -3863 16081 -3811
rect 14423 -4171 14475 -3911
rect 14481 -4271 16081 -4219
rect 16066 -4389 16206 -4337
rect 14193 -5219 14333 -5141
rect 16231 -5220 16370 -5141
<< metal2 >>
rect 13457 1921 15921 1931
rect 13614 1918 15921 1921
rect 13614 1861 14296 1918
rect 15896 1861 15921 1918
rect 13457 1851 15921 1861
rect 13386 1813 14290 1823
rect 2205 1796 2425 1806
rect 2205 1598 2425 1608
rect 5688 1796 5908 1806
rect 5688 1598 5908 1608
rect 9176 1796 9396 1806
rect 9176 1598 9396 1608
rect 13386 1804 14238 1813
rect 13386 1616 13404 1804
rect 13624 1616 14238 1804
rect 13386 1613 14238 1616
rect 13386 1603 14290 1613
rect 15900 1813 15966 1823
rect 15956 1613 15966 1813
rect 15900 1603 15966 1613
rect 13457 1565 15921 1575
rect 13614 1508 14296 1565
rect 15896 1508 15921 1565
rect 13614 1505 15921 1508
rect 13457 1495 15921 1505
rect 13457 1389 15916 1399
rect 13614 1386 15916 1389
rect 13614 1329 14296 1386
rect 15896 1329 15916 1386
rect 13457 1319 15916 1329
rect 13447 1033 15916 1043
rect 13447 976 13457 1033
rect 5504 973 13457 976
rect 13614 976 14297 1033
rect 15897 976 15916 1033
rect 13614 973 15916 976
rect 5504 966 15916 973
rect 5661 906 12471 966
rect 12628 963 15916 966
rect 12628 906 13624 963
rect 5504 896 13624 906
rect 13447 867 13624 896
rect 2349 857 13377 867
rect 2349 853 13220 857
rect 5549 797 5835 853
rect 9035 797 9321 853
rect 12521 797 13220 853
rect 2349 787 13377 797
rect 13447 857 15916 867
rect 13447 797 13457 857
rect 13614 854 15916 857
rect 13614 797 14296 854
rect 15896 797 15916 854
rect 13447 788 15916 797
rect 13457 787 15916 788
rect 2289 749 2345 759
rect 2289 539 2345 549
rect 5553 749 5609 759
rect 5553 539 5609 549
rect 5775 749 5831 759
rect 5775 539 5831 549
rect 9261 749 9317 759
rect 9261 539 9317 549
rect 12525 749 12581 759
rect 12525 539 12581 549
rect 2349 501 13377 511
rect 5549 445 5835 501
rect 9035 445 9321 501
rect 12521 445 13220 501
rect 2349 441 13220 445
rect 2349 431 13377 441
rect 13457 501 15916 511
rect 13614 444 14296 501
rect 15896 444 15916 501
rect 13614 441 15916 444
rect 13457 431 15916 441
rect 2349 325 13377 335
rect 2349 321 13220 325
rect 5549 265 5835 321
rect 9035 265 9321 321
rect 12521 265 13220 321
rect 2349 255 13377 265
rect 13457 325 15921 335
rect 13614 322 15921 325
rect 13614 265 14296 322
rect 15896 265 15921 322
rect 13457 255 15921 265
rect 5553 217 5609 227
rect 5553 7 5609 17
rect 12525 217 12581 227
rect 12525 7 12581 17
rect 15900 217 15966 227
rect 15956 17 15966 217
rect 15900 7 15966 17
rect 2349 -31 13377 -21
rect 5549 -87 5835 -31
rect 9035 -87 9321 -31
rect 12521 -87 13220 -31
rect 2349 -91 13220 -87
rect 2349 -101 13377 -91
rect 13457 -31 15924 -21
rect 13614 -88 14296 -31
rect 15896 -88 15924 -31
rect 13614 -91 15924 -88
rect 13457 -101 15924 -91
rect 5504 -139 13614 -129
rect 5661 -199 12471 -139
rect 12628 -199 13457 -139
rect 5504 -209 13614 -199
rect 7668 -765 16007 -755
rect 7668 -821 7678 -765
rect 7818 -821 13229 -765
rect 13369 -821 15857 -765
rect 15997 -821 16007 -765
rect 7668 -831 16007 -821
rect 8554 -903 13624 -894
rect 8554 -959 8565 -903
rect 8705 -904 13624 -903
rect 8705 -959 12229 -904
rect 8554 -960 12229 -959
rect 12369 -905 13624 -904
rect 12369 -960 13467 -905
rect 8554 -961 13467 -960
rect 13607 -961 13624 -905
rect 8554 -970 13624 -961
rect 7074 -1103 9806 -1093
rect 7074 -1107 8842 -1103
rect 7674 -1159 7960 -1107
rect 8560 -1159 8842 -1107
rect 8982 -1107 9806 -1103
rect 8982 -1159 9206 -1107
rect 7074 -1169 9806 -1159
rect 10452 -1105 12379 -1097
rect 10452 -1107 12229 -1105
rect 12052 -1159 12229 -1107
rect 10452 -1161 12229 -1159
rect 12369 -1161 12379 -1105
rect 10452 -1169 12379 -1161
rect 12808 -1106 13387 -1099
rect 12808 -1107 13228 -1106
rect 13008 -1159 13228 -1107
rect 12808 -1162 13228 -1159
rect 13368 -1162 13387 -1106
rect 12808 -1169 13387 -1162
rect 7678 -1207 7734 -1197
rect 7678 -1417 7734 -1407
rect 8564 -1207 8620 -1197
rect 8564 -1417 8620 -1407
rect 12058 -1207 12110 -1197
rect 12110 -1279 12599 -1269
rect 12110 -1335 12449 -1279
rect 12589 -1335 12599 -1279
rect 12110 -1345 12599 -1335
rect 12058 -1417 12110 -1407
rect 7074 -1455 9806 -1445
rect 7674 -1507 7960 -1455
rect 8560 -1507 8842 -1455
rect 7074 -1511 8842 -1507
rect 8982 -1507 9206 -1455
rect 8982 -1511 9806 -1507
rect 7074 -1521 9806 -1511
rect 10452 -1455 12379 -1445
rect 12052 -1507 12226 -1455
rect 10452 -1511 12226 -1507
rect 12366 -1511 12379 -1455
rect 10452 -1517 12379 -1511
rect 13447 -1750 14579 -1740
rect 8835 -1816 9808 -1806
rect 8835 -1872 8842 -1816
rect 8982 -1820 9808 -1816
rect 13447 -1810 13457 -1750
rect 13614 -1810 14421 -1750
rect 14578 -1810 14579 -1750
rect 13447 -1820 14579 -1810
rect 8982 -1872 9212 -1820
rect 8835 -1882 9808 -1872
rect 10452 -1856 12599 -1846
rect 10452 -1860 12449 -1856
rect 9148 -1920 9204 -1910
rect 12052 -1912 12449 -1860
rect 12589 -1912 12599 -1856
rect 10452 -1922 12599 -1912
rect 12808 -1853 13387 -1845
rect 12808 -1855 13228 -1853
rect 13008 -1907 13228 -1855
rect 12808 -1909 13228 -1907
rect 13368 -1909 13387 -1853
rect 14183 -1863 14340 -1859
rect 12808 -1917 13387 -1909
rect 14177 -1869 16081 -1863
rect 14177 -1929 14183 -1869
rect 14340 -1873 16081 -1869
rect 14340 -1925 14481 -1873
rect 14340 -1929 16081 -1925
rect 14177 -1935 16081 -1929
rect 14183 -1939 14340 -1935
rect 9148 -2130 9204 -2120
rect 10392 -1960 10448 -1950
rect 8628 -2168 9804 -2158
rect 8628 -2224 8656 -2168
rect 8983 -2220 9208 -2168
rect 10392 -2170 10448 -2160
rect 14421 -1973 14477 -1963
rect 8983 -2224 9804 -2220
rect 8628 -2234 9804 -2224
rect 10452 -2207 13008 -2198
rect 10452 -2208 12449 -2207
rect 12052 -2260 12449 -2208
rect 10452 -2263 12449 -2260
rect 12589 -2208 13008 -2207
rect 12589 -2260 12808 -2208
rect 14421 -2243 14477 -2233
rect 12589 -2263 13008 -2260
rect 10452 -2270 13008 -2263
rect 14183 -2271 14340 -2267
rect 14177 -2277 16081 -2271
rect 12750 -2308 12802 -2298
rect 11236 -2400 12750 -2390
rect 11376 -2456 12750 -2400
rect 11236 -2466 12750 -2456
rect 8408 -2582 11938 -2572
rect 8408 -2638 8418 -2582
rect 8558 -2638 9064 -2582
rect 9204 -2586 11938 -2582
rect 9204 -2638 9566 -2586
rect 10166 -2638 10452 -2586
rect 11052 -2638 11338 -2586
rect 8408 -2648 11938 -2638
rect 9506 -2686 9562 -2676
rect 9506 -2896 9562 -2886
rect 10392 -2686 10448 -2676
rect 10392 -2896 10448 -2886
rect 11278 -2686 11334 -2676
rect 11278 -2896 11334 -2886
rect 14177 -2337 14183 -2277
rect 14340 -2281 16081 -2277
rect 14340 -2333 14481 -2281
rect 14340 -2337 16081 -2333
rect 14177 -2343 16081 -2337
rect 14183 -2347 14340 -2343
rect 13210 -2396 14578 -2386
rect 13210 -2456 13220 -2396
rect 13377 -2456 14421 -2396
rect 13210 -2466 14578 -2456
rect 16221 -2509 16378 -2505
rect 14481 -2515 16385 -2509
rect 14481 -2519 16221 -2515
rect 16081 -2571 16221 -2519
rect 14481 -2575 16221 -2571
rect 16378 -2575 16385 -2515
rect 14481 -2581 16385 -2575
rect 16221 -2585 16378 -2581
rect 14421 -2619 14477 -2609
rect 14421 -2889 14477 -2879
rect 12750 -2918 12802 -2908
rect 16221 -2917 16378 -2913
rect 14481 -2923 16385 -2917
rect 9054 -2934 11938 -2924
rect 9054 -2990 9064 -2934
rect 9204 -2986 9566 -2934
rect 10166 -2986 10452 -2934
rect 11052 -2986 11338 -2934
rect 14481 -2927 16221 -2923
rect 9204 -2990 11938 -2986
rect 9054 -3000 11938 -2990
rect 12439 -2952 13008 -2946
rect 12439 -3008 12448 -2952
rect 12588 -2956 13008 -2952
rect 12588 -3008 12808 -2956
rect 16081 -2979 16221 -2927
rect 14481 -2983 16221 -2979
rect 16378 -2983 16385 -2923
rect 14481 -2989 16385 -2983
rect 16221 -2993 16378 -2989
rect 12439 -3017 13008 -3008
rect 13210 -3042 14578 -3032
rect 13210 -3102 13220 -3042
rect 13377 -3102 14421 -3042
rect 13210 -3112 14578 -3102
rect 8865 -3139 9572 -3129
rect 8865 -3199 8875 -3139
rect 9032 -3199 9405 -3139
rect 9562 -3199 9572 -3139
rect 16221 -3155 16378 -3151
rect 8865 -3209 9572 -3199
rect 14481 -3161 16385 -3155
rect 14481 -3165 16221 -3161
rect 16081 -3217 16221 -3165
rect 14481 -3221 16221 -3217
rect 16378 -3221 16385 -3161
rect 14481 -3227 16385 -3221
rect 16221 -3231 16378 -3227
rect 14421 -3265 14477 -3255
rect 8865 -3368 13208 -3362
rect 8865 -3428 8875 -3368
rect 9032 -3372 13208 -3368
rect 9032 -3424 9208 -3372
rect 9032 -3428 13208 -3424
rect 8865 -3434 13208 -3428
rect 9150 -3472 9202 -3462
rect 14421 -3535 14477 -3525
rect 16221 -3563 16378 -3559
rect 14481 -3569 16385 -3563
rect 14481 -3573 16221 -3569
rect 16081 -3625 16221 -3573
rect 14481 -3628 16221 -3625
rect 16378 -3628 16385 -3569
rect 14481 -3635 16385 -3628
rect 16221 -3639 16378 -3635
rect 9150 -3682 9202 -3672
rect 13447 -3688 14578 -3678
rect 8483 -3716 13208 -3710
rect 8483 -3776 8875 -3716
rect 9032 -3720 13208 -3716
rect 9032 -3772 9208 -3720
rect 13447 -3748 13457 -3688
rect 13614 -3748 14421 -3688
rect 13447 -3758 14578 -3748
rect 9032 -3776 13208 -3772
rect 8483 -3786 13208 -3776
rect 14183 -3801 14340 -3798
rect 14177 -3808 16081 -3801
rect 14177 -3868 14183 -3808
rect 14340 -3811 16081 -3808
rect 14340 -3863 14481 -3811
rect 14340 -3868 16081 -3863
rect 14177 -3873 16081 -3868
rect 8865 -3882 13208 -3876
rect 14183 -3878 14340 -3873
rect 7385 -3926 8805 -3917
rect 7385 -3986 8639 -3926
rect 8796 -3986 8805 -3926
rect 8865 -3942 8875 -3882
rect 9032 -3886 13208 -3882
rect 9032 -3938 9208 -3886
rect 9032 -3942 13208 -3938
rect 8865 -3948 13208 -3942
rect 14421 -3911 14477 -3901
rect 7385 -3993 8805 -3986
rect 9148 -3986 9204 -3976
rect 14421 -4181 14477 -4171
rect 9148 -4196 9204 -4186
rect 6953 -4211 7031 -4201
rect 14183 -4209 14340 -4205
rect 14183 -4215 16081 -4209
rect 8865 -4230 13208 -4224
rect 7031 -4345 7157 -4269
rect 8865 -4290 8875 -4230
rect 9032 -4234 13208 -4230
rect 9032 -4286 9208 -4234
rect 14340 -4219 16081 -4215
rect 14340 -4271 14481 -4219
rect 14340 -4275 16081 -4271
rect 14183 -4281 16081 -4275
rect 14183 -4285 14340 -4281
rect 9032 -4290 13208 -4286
rect 8865 -4296 13208 -4290
rect 9104 -4334 16206 -4324
rect 6953 -4361 7031 -4351
rect 9244 -4337 16206 -4334
rect 9244 -4389 16066 -4337
rect 9244 -4390 16206 -4389
rect 9104 -4400 16206 -4390
rect 14193 -5141 14333 -5131
rect 14193 -5229 14333 -5219
rect 16231 -5141 16370 -5131
rect 16231 -5230 16370 -5220
<< via2 >>
rect 13457 1861 13614 1921
rect 2205 1608 2425 1796
rect 5688 1608 5908 1796
rect 9176 1608 9396 1796
rect 15900 1613 15902 1813
rect 15902 1613 15954 1813
rect 15954 1613 15956 1813
rect 13457 1505 13614 1565
rect 13457 1329 13614 1389
rect 13457 973 13614 1033
rect 5504 906 5661 966
rect 12471 906 12628 966
rect 13220 797 13377 857
rect 13457 797 13614 857
rect 2289 549 2291 749
rect 2291 549 2343 749
rect 2343 549 2345 749
rect 5553 549 5555 749
rect 5555 549 5607 749
rect 5607 549 5609 749
rect 5775 549 5777 749
rect 5777 549 5829 749
rect 5829 549 5831 749
rect 9261 549 9263 749
rect 9263 549 9315 749
rect 9315 549 9317 749
rect 12525 549 12527 749
rect 12527 549 12579 749
rect 12579 549 12581 749
rect 13220 441 13377 501
rect 13457 441 13614 501
rect 13220 265 13377 325
rect 13457 265 13614 325
rect 5553 17 5555 217
rect 5555 17 5607 217
rect 5607 17 5609 217
rect 12525 17 12527 217
rect 12527 17 12579 217
rect 12579 17 12581 217
rect 15900 17 15902 217
rect 15902 17 15954 217
rect 15954 17 15956 217
rect 13220 -91 13377 -31
rect 13457 -91 13614 -31
rect 5504 -199 5661 -139
rect 12471 -199 12628 -139
rect 13457 -199 13614 -139
rect 7678 -821 7818 -765
rect 13229 -821 13369 -765
rect 15857 -821 15997 -765
rect 8565 -959 8705 -903
rect 12229 -960 12369 -904
rect 13467 -961 13607 -905
rect 8842 -1159 8982 -1103
rect 12229 -1161 12369 -1105
rect 13228 -1162 13368 -1106
rect 7678 -1407 7680 -1207
rect 7680 -1407 7732 -1207
rect 7732 -1407 7734 -1207
rect 8564 -1407 8566 -1207
rect 8566 -1407 8618 -1207
rect 8618 -1407 8620 -1207
rect 12449 -1335 12589 -1279
rect 8842 -1511 8982 -1455
rect 12226 -1511 12366 -1455
rect 8842 -1872 8982 -1816
rect 13457 -1810 13614 -1750
rect 14421 -1810 14578 -1750
rect 9148 -2120 9150 -1920
rect 9150 -2120 9202 -1920
rect 9202 -2120 9204 -1920
rect 12449 -1912 12589 -1856
rect 13228 -1909 13368 -1853
rect 14183 -1929 14340 -1869
rect 8656 -2224 8983 -2168
rect 10392 -2160 10394 -1960
rect 10394 -2160 10446 -1960
rect 10446 -2160 10448 -1960
rect 12449 -2263 12589 -2207
rect 14421 -2233 14423 -1973
rect 14423 -2233 14475 -1973
rect 14475 -2233 14477 -1973
rect 11236 -2456 11376 -2400
rect 8418 -2638 8558 -2582
rect 9064 -2638 9204 -2582
rect 9506 -2886 9508 -2686
rect 9508 -2886 9560 -2686
rect 9560 -2886 9562 -2686
rect 10392 -2886 10394 -2686
rect 10394 -2886 10446 -2686
rect 10446 -2886 10448 -2686
rect 11278 -2886 11280 -2686
rect 11280 -2886 11332 -2686
rect 11332 -2886 11334 -2686
rect 14183 -2337 14340 -2277
rect 13220 -2456 13377 -2396
rect 14421 -2456 14578 -2396
rect 16221 -2575 16378 -2515
rect 14421 -2879 14423 -2619
rect 14423 -2879 14475 -2619
rect 14475 -2879 14477 -2619
rect 9064 -2990 9204 -2934
rect 12448 -3008 12588 -2952
rect 16221 -2983 16378 -2923
rect 13220 -3102 13377 -3042
rect 14421 -3102 14578 -3042
rect 8875 -3199 9032 -3139
rect 9405 -3199 9562 -3139
rect 16221 -3221 16378 -3161
rect 8875 -3428 9032 -3368
rect 14421 -3525 14423 -3265
rect 14423 -3525 14475 -3265
rect 14475 -3525 14477 -3265
rect 16221 -3628 16378 -3569
rect 8875 -3776 9032 -3716
rect 13457 -3748 13614 -3688
rect 14421 -3748 14578 -3688
rect 14183 -3868 14340 -3808
rect 8639 -3986 8796 -3926
rect 8875 -3942 9032 -3882
rect 9148 -4186 9150 -3986
rect 9150 -4186 9202 -3986
rect 9202 -4186 9204 -3986
rect 14421 -4171 14423 -3911
rect 14423 -4171 14475 -3911
rect 14475 -4171 14477 -3911
rect 8875 -4290 9032 -4230
rect 14183 -4275 14340 -4215
rect 9104 -4390 9244 -4334
rect 14193 -5219 14333 -5141
rect 16231 -5220 16370 -5141
<< metal3 >>
rect 13447 1921 13624 1932
rect 13447 1861 13457 1921
rect 13614 1861 13624 1921
rect 2195 1796 2435 1801
rect 2195 1608 2205 1796
rect 2425 1608 2435 1796
rect 2195 1603 2435 1608
rect 5678 1796 5918 1801
rect 5678 1608 5688 1796
rect 5908 1608 5918 1796
rect 5678 1603 5918 1608
rect 9166 1796 9406 1801
rect 9166 1608 9176 1796
rect 9396 1608 9406 1796
rect 9166 1603 9406 1608
rect 2279 749 2355 1603
rect 5494 966 5671 971
rect 5494 906 5504 966
rect 5661 906 5671 966
rect 5494 901 5671 906
rect 2279 549 2289 749
rect 2345 549 2355 749
rect 2279 544 2355 549
rect 5543 749 5619 901
rect 5543 549 5553 749
rect 5609 549 5619 749
rect 5543 217 5619 549
rect 5765 749 5841 1603
rect 5765 549 5775 749
rect 5831 549 5841 749
rect 5765 544 5841 549
rect 9251 749 9327 1603
rect 13447 1565 13624 1861
rect 13447 1505 13457 1565
rect 13614 1505 13624 1565
rect 13447 1389 13624 1505
rect 13447 1329 13457 1389
rect 13614 1329 13624 1389
rect 13447 1033 13624 1329
rect 13447 973 13457 1033
rect 13614 973 13624 1033
rect 12461 966 12638 971
rect 12461 906 12471 966
rect 12628 906 12638 966
rect 12461 901 12638 906
rect 9251 549 9261 749
rect 9317 549 9327 749
rect 9251 544 9327 549
rect 12515 749 12591 901
rect 12515 549 12525 749
rect 12581 549 12591 749
rect 5543 17 5553 217
rect 5609 17 5619 217
rect 5543 -134 5619 17
rect 12515 217 12591 549
rect 12515 17 12525 217
rect 12581 17 12591 217
rect 12515 -134 12591 17
rect 13210 857 13387 868
rect 13210 797 13220 857
rect 13377 797 13387 857
rect 13210 501 13387 797
rect 13210 441 13220 501
rect 13377 441 13387 501
rect 13210 325 13387 441
rect 13210 265 13220 325
rect 13377 265 13387 325
rect 13210 -31 13387 265
rect 13210 -91 13220 -31
rect 13377 -91 13387 -31
rect 5494 -139 5671 -134
rect 5494 -199 5504 -139
rect 5661 -199 5671 -139
rect 5494 -204 5671 -199
rect 12461 -139 12638 -134
rect 12461 -199 12471 -139
rect 12628 -199 12638 -139
rect 12461 -204 12638 -199
rect 7668 -765 7828 -755
rect 7668 -821 7678 -765
rect 7818 -821 7828 -765
rect 7668 -1207 7828 -821
rect 13210 -765 13387 -91
rect 13210 -821 13229 -765
rect 13369 -821 13387 -765
rect 7668 -1407 7678 -1207
rect 7734 -1407 7828 -1207
rect 7668 -1412 7828 -1407
rect 8554 -903 8714 -894
rect 8554 -959 8565 -903
rect 8705 -959 8714 -903
rect 8554 -1207 8714 -959
rect 12219 -904 12379 -894
rect 12219 -960 12229 -904
rect 12369 -960 12379 -904
rect 8554 -1407 8564 -1207
rect 8620 -1407 8714 -1207
rect 8554 -1412 8714 -1407
rect 8832 -1103 8992 -1093
rect 8832 -1159 8842 -1103
rect 8982 -1159 8992 -1103
rect 8832 -1455 8992 -1159
rect 8832 -1511 8842 -1455
rect 8982 -1511 8992 -1455
rect 8832 -1816 8992 -1511
rect 12219 -1105 12379 -960
rect 12219 -1161 12229 -1105
rect 12369 -1161 12379 -1105
rect 12219 -1455 12379 -1161
rect 13210 -1106 13387 -821
rect 13210 -1162 13228 -1106
rect 13368 -1162 13387 -1106
rect 12219 -1511 12226 -1455
rect 12366 -1511 12379 -1455
rect 12219 -1517 12379 -1511
rect 12439 -1279 12599 -1269
rect 12439 -1335 12449 -1279
rect 12589 -1335 12599 -1279
rect 8832 -1872 8842 -1816
rect 8982 -1872 8992 -1816
rect 8832 -2158 8992 -1872
rect 12439 -1856 12599 -1335
rect 12439 -1912 12449 -1856
rect 12589 -1912 12599 -1856
rect 8628 -2168 8992 -2158
rect 8628 -2224 8656 -2168
rect 8983 -2224 8992 -2168
rect 8628 -2234 8992 -2224
rect 9054 -1920 9214 -1915
rect 9054 -2120 9148 -1920
rect 9204 -2120 9214 -1920
rect 8408 -2582 8568 -2577
rect 8408 -2638 8418 -2582
rect 8558 -2638 8568 -2582
rect 8408 -2643 8568 -2638
rect 8628 -3926 8805 -2234
rect 9054 -2582 9214 -2120
rect 9054 -2638 9064 -2582
rect 9204 -2638 9214 -2582
rect 9054 -2934 9214 -2638
rect 10382 -1960 10458 -1955
rect 10382 -2160 10392 -1960
rect 10448 -2160 10458 -1960
rect 9054 -2990 9064 -2934
rect 9204 -2990 9214 -2934
rect 9054 -2996 9214 -2990
rect 9395 -2681 9509 -2680
rect 9395 -2686 9572 -2681
rect 9395 -2886 9506 -2686
rect 9562 -2886 9572 -2686
rect 8628 -3986 8639 -3926
rect 8796 -3986 8805 -3926
rect 8628 -3993 8805 -3986
rect 8865 -3139 9042 -3129
rect 8865 -3199 8875 -3139
rect 9032 -3199 9042 -3139
rect 8865 -3368 9042 -3199
rect 9395 -3139 9572 -2886
rect 10382 -2686 10458 -2160
rect 12439 -2207 12599 -1912
rect 12439 -2263 12449 -2207
rect 12589 -2263 12599 -2207
rect 11226 -2400 11386 -2395
rect 11226 -2456 11236 -2400
rect 11376 -2456 11386 -2400
rect 11226 -2461 11386 -2456
rect 10382 -2886 10392 -2686
rect 10448 -2886 10458 -2686
rect 10382 -2891 10458 -2886
rect 11268 -2686 11344 -2461
rect 11268 -2886 11278 -2686
rect 11334 -2886 11344 -2686
rect 11268 -2891 11344 -2886
rect 12439 -2952 12599 -2263
rect 12439 -3008 12448 -2952
rect 12588 -3008 12599 -2952
rect 12439 -3017 12599 -3008
rect 13210 -1853 13387 -1162
rect 13210 -1909 13228 -1853
rect 13368 -1909 13387 -1853
rect 13210 -2396 13387 -1909
rect 13210 -2456 13220 -2396
rect 13377 -2456 13387 -2396
rect 13210 -3042 13387 -2456
rect 13210 -3102 13220 -3042
rect 13377 -3102 13387 -3042
rect 13210 -3112 13387 -3102
rect 13447 857 13624 973
rect 13447 797 13457 857
rect 13614 797 13624 857
rect 13447 501 13624 797
rect 13447 441 13457 501
rect 13614 441 13624 501
rect 13447 325 13624 441
rect 13447 265 13457 325
rect 13614 265 13624 325
rect 13447 -31 13624 265
rect 13447 -91 13457 -31
rect 13614 -91 13624 -31
rect 13447 -139 13624 -91
rect 13447 -199 13457 -139
rect 13614 -199 13624 -139
rect 13447 -905 13624 -199
rect 15890 1813 15966 1818
rect 15890 1613 15900 1813
rect 15956 1613 15966 1813
rect 15890 217 15966 1613
rect 15890 17 15900 217
rect 15956 17 15966 217
rect 15890 -760 15966 17
rect 15847 -765 16007 -760
rect 15847 -821 15857 -765
rect 15997 -821 16007 -765
rect 15847 -831 16007 -821
rect 13447 -961 13467 -905
rect 13607 -961 13624 -905
rect 13447 -1750 13624 -961
rect 13447 -1810 13457 -1750
rect 13614 -1810 13624 -1750
rect 9395 -3199 9405 -3139
rect 9562 -3199 9572 -3139
rect 9395 -3209 9572 -3199
rect 8865 -3428 8875 -3368
rect 9032 -3428 9042 -3368
rect 8865 -3716 9042 -3428
rect 8865 -3776 8875 -3716
rect 9032 -3776 9042 -3716
rect 13447 -3688 13624 -1810
rect 14411 -1750 14588 -1745
rect 14411 -1810 14421 -1750
rect 14578 -1810 14588 -1750
rect 14411 -1815 14588 -1810
rect 13447 -3748 13457 -3688
rect 13614 -3748 13624 -3688
rect 13447 -3758 13624 -3748
rect 14173 -1869 14350 -1864
rect 14173 -1929 14183 -1869
rect 14340 -1929 14350 -1869
rect 14173 -2277 14350 -1929
rect 14411 -1973 14487 -1815
rect 14411 -2233 14421 -1973
rect 14477 -2233 14487 -1973
rect 14411 -2238 14487 -2233
rect 14173 -2337 14183 -2277
rect 14340 -2337 14350 -2277
rect 8865 -3882 9042 -3776
rect 8865 -3942 8875 -3882
rect 9032 -3942 9042 -3882
rect 8865 -4230 9042 -3942
rect 14173 -3808 14350 -2337
rect 14411 -2391 14487 -2390
rect 14411 -2396 14588 -2391
rect 14411 -2456 14421 -2396
rect 14578 -2456 14588 -2396
rect 14411 -2461 14588 -2456
rect 14411 -2619 14487 -2461
rect 14411 -2879 14421 -2619
rect 14477 -2879 14487 -2619
rect 14411 -2884 14487 -2879
rect 16211 -2515 16388 -2510
rect 16211 -2575 16221 -2515
rect 16378 -2575 16388 -2515
rect 16211 -2923 16388 -2575
rect 16211 -2983 16221 -2923
rect 16378 -2983 16388 -2923
rect 14411 -3042 14588 -3037
rect 14411 -3102 14421 -3042
rect 14578 -3102 14588 -3042
rect 14411 -3107 14588 -3102
rect 14411 -3265 14487 -3107
rect 14411 -3525 14421 -3265
rect 14477 -3525 14487 -3265
rect 14411 -3531 14487 -3525
rect 16211 -3161 16388 -2983
rect 16211 -3221 16221 -3161
rect 16378 -3221 16388 -3161
rect 16211 -3569 16388 -3221
rect 16211 -3628 16221 -3569
rect 16378 -3628 16388 -3569
rect 14173 -3868 14183 -3808
rect 14340 -3868 14350 -3808
rect 8865 -4290 8875 -4230
rect 9032 -4290 9042 -4230
rect 8865 -4296 9042 -4290
rect 9138 -3986 9214 -3981
rect 9138 -4186 9148 -3986
rect 9204 -4186 9214 -3986
rect 9138 -4329 9214 -4186
rect 14173 -4215 14350 -3868
rect 14411 -3688 14588 -3683
rect 14411 -3748 14421 -3688
rect 14578 -3748 14588 -3688
rect 14411 -3753 14588 -3748
rect 14411 -3911 14487 -3753
rect 14411 -4171 14421 -3911
rect 14477 -4171 14487 -3911
rect 14411 -4176 14487 -4171
rect 14173 -4275 14183 -4215
rect 14340 -4275 14350 -4215
rect 9094 -4334 9254 -4329
rect 9094 -4390 9104 -4334
rect 9244 -4390 9254 -4334
rect 9094 -4395 9254 -4390
rect 14173 -5141 14350 -4275
rect 14173 -5219 14193 -5141
rect 14333 -5219 14350 -5141
rect 14173 -5229 14350 -5219
rect 16211 -5141 16388 -3628
rect 16211 -5220 16231 -5141
rect 16370 -5220 16388 -5141
rect 16211 -5230 16388 -5220
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  D1
timestamp 1712928760
transform 0 1 14263 -1 0 -5180
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  D3
timestamp 1712928760
transform 1 0 6992 0 1 -4281
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0
timestamp 1712928760
transform 0 1 16300 -1 0 -5180
box -183 -208 183 208
use trans_gate  x1
timestamp 1712947935
transform 1 0 5910 0 1 -2437
box 1220 -2096 2736 522
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[0]
timestamp 1712777902
transform 1 0 15281 0 1 -2103
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[1]
timestamp 1712777902
transform 1 0 15281 0 1 -4041
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[0]
timestamp 1712777902
transform 1 0 15281 0 1 -2749
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[1]
timestamp 1712777902
transform 1 0 15281 0 1 -3395
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[0]
timestamp 1712777902
transform 1 0 15096 0 1 1181
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[1]
timestamp 1712777902
transform 1 0 15096 0 1 649
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM4[0]
timestamp 1712777902
transform 1 0 7435 0 1 649
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1712777902
transform 1 0 7435 0 1 117
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[0]
timestamp 1712777902
transform 1 0 15096 0 1 1713
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[1]
timestamp 1712777902
transform 1 0 15096 0 1 117
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[0]
timestamp 1712777902
transform 1 0 3949 0 1 649
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1712777902
transform 1 0 3949 0 1 117
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[2]
timestamp 1712777902
transform 1 0 10921 0 1 649
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1712777902
transform 1 0 10921 0 1 117
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1712777902
transform 1 0 11252 0 1 -1307
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_697RXD  XM8
timestamp 1712777902
transform 1 0 11252 0 1 -2060
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1712777902
transform 1 0 12908 0 1 -1507
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1712777902
transform 1 0 12908 0 1 -2608
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1712777902
transform 1 0 11208 0 1 -3572
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1712777902
transform 1 0 11208 0 1 -4086
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1712847059
transform 1 0 9858 0 1 -2786
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1712847059
transform 1 0 10744 0 1 -2786
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1712856153
transform 1 0 8260 0 1 -1307
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1712856153
transform 1 0 7374 0 1 -1307
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1712847059
transform 1 0 11630 0 1 -2786
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1712856153
transform 1 0 9506 0 1 -1307
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1712847059
transform 1 0 9508 0 1 -2020
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[0]
timestamp 1712777902
transform 1 0 13910 0 1 2245
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[1]
timestamp 1712777902
transform 1 0 13910 0 1 1713
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[2]
timestamp 1712777902
transform 1 0 13910 0 1 1181
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[3]
timestamp 1712777902
transform 1 0 13910 0 1 649
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712777902
transform 1 0 13910 0 1 117
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712777902
transform 1 0 13910 0 1 -415
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712777902
transform 1 0 16282 0 1 2245
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712777902
transform 1 0 16282 0 1 1713
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712777902
transform 1 0 16282 0 1 1181
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712777902
transform 1 0 16282 0 1 649
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712777902
transform 1 0 16282 0 1 117
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712777902
transform 1 0 16282 0 1 -415
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712777902
transform 1 0 1963 0 1 1181
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712777902
transform 1 0 1963 0 1 649
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712777902
transform 1 0 1963 0 1 117
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712777902
transform 1 0 1963 0 1 -415
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[16]
timestamp 1712777902
transform 1 0 12907 0 1 1181
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[17]
timestamp 1712777902
transform 1 0 12907 0 1 649
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[18]
timestamp 1712777902
transform 1 0 12907 0 1 117
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[19]
timestamp 1712777902
transform 1 0 12907 0 1 -415
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[0]
timestamp 1712777902
transform 1 0 15096 0 1 2245
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[1]
timestamp 1712777902
transform 1 0 15096 0 1 -415
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712777902
transform 1 0 3949 0 1 1181
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712777902
transform 1 0 7435 0 1 1181
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712777902
transform 1 0 10921 0 1 1181
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712777902
transform 1 0 3949 0 1 -415
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712777902
transform 1 0 7435 0 1 -415
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712777902
transform 1 0 10921 0 1 -415
box -1796 -319 1796 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712777902
transform 1 0 13943 0 1 -1487
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712777902
transform 1 0 13943 0 1 -4657
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712777902
transform 1 0 16619 0 1 -1487
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712777902
transform 1 0 16619 0 1 -4657
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712777902
transform 1 0 15281 0 1 -1487
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712777902
transform 1 0 15281 0 1 -4657
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712777902
transform 1 0 13943 0 1 -2103
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712777902
transform 1 0 13943 0 1 -2749
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712777902
transform 1 0 13943 0 1 -3395
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712777902
transform 1 0 13943 0 1 -4041
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[4]
timestamp 1712777902
transform 1 0 16619 0 1 -2103
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[5]
timestamp 1712777902
transform 1 0 16619 0 1 -2749
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[6]
timestamp 1712777902
transform 1 0 16619 0 1 -3395
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[7]
timestamp 1712777902
transform 1 0 16619 0 1 -4041
box -328 -388 328 388
<< labels >>
flabel metal1 7108 -3786 7157 -3710 0 FreeSans 1280 0 0 0 ibias
port 6 nsew
flabel metal3 14173 -5229 14350 -5131 0 FreeSans 1280 0 0 0 vref
port 3 nsew
flabel metal3 16211 -5230 16388 -5131 0 FreeSans 1280 0 0 0 vin
port 4 nsew
flabel metal2 6953 -4361 7031 -4201 0 FreeSans 1280 0 0 0 ena
port 5 nsew
flabel metal1 6845 -5327 7446 -4931 0 FreeSans 1600 0 0 0 vss
port 7 nsew
flabel metal1 1703 2134 2208 2528 0 FreeSans 1600 0 0 0 dvdd
port 1 nsew
flabel metal1 16272 -1017 16661 -839 0 FreeSans 1600 0 0 0 out
port 8 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712752659
<< nwell >>
rect 15899 1675 15954 1683
rect 14281 1437 15936 1444
rect 15918 1365 15936 1437
<< metal1 >>
rect 13758 2246 16434 2292
rect 13758 1964 13804 2246
rect 14016 1964 14062 2246
rect 14190 1964 14290 2246
rect 15902 1964 15948 2246
rect 16130 1964 16176 2246
rect 16388 1964 16434 2246
rect 13758 1918 16434 1964
rect 13758 1760 13804 1918
rect 14016 1760 14062 1918
rect 13758 1714 13822 1760
rect 14001 1714 14062 1760
rect 13758 1432 13804 1714
rect 14016 1432 14062 1714
rect 13758 1386 13826 1432
rect 14004 1386 14062 1432
rect 13758 1228 13804 1386
rect 14016 1228 14062 1386
rect 1811 1182 13059 1228
rect 1811 900 1857 1182
rect 2069 900 2115 1182
rect 2265 900 2343 1182
rect 5555 900 5601 1182
rect 5751 900 5829 1182
rect 9041 900 9087 1182
rect 9237 900 9315 1182
rect 12527 900 12573 1182
rect 12755 900 12801 1182
rect 13013 900 13059 1182
rect 1811 854 13059 900
rect 1811 696 1857 854
rect 2069 696 2115 854
rect 1811 650 1888 696
rect 2051 650 2115 696
rect 1811 368 1857 650
rect 2069 368 2115 650
rect 1811 322 1884 368
rect 2053 322 2115 368
rect 1811 164 1857 322
rect 2069 164 2115 322
rect 1811 118 1885 164
rect 2056 118 2115 164
rect 1811 -164 1857 118
rect 2069 -164 2115 118
rect 1811 -210 1889 -164
rect 2052 -210 2115 -164
rect 1811 -368 1857 -210
rect 2069 -368 2115 -210
rect 2265 -368 2311 854
rect 2339 657 2349 713
rect 5549 657 5559 713
rect 2339 650 5559 657
rect 5545 409 5555 609
rect 5607 409 5617 609
rect 2339 361 5559 368
rect 2339 305 2349 361
rect 5549 305 5559 361
rect 2339 125 2349 181
rect 5549 125 5559 181
rect 2339 118 5559 125
rect 5545 -123 5555 77
rect 5607 -123 5617 77
rect 2339 -171 5559 -164
rect 2339 -227 2349 -171
rect 5549 -227 5559 -171
rect 5751 -368 5797 854
rect 5825 657 5835 713
rect 9035 657 9087 713
rect 5825 650 9087 657
rect 9041 609 9087 650
rect 9041 368 9087 409
rect 5825 361 9087 368
rect 5825 305 5835 361
rect 9035 305 9087 361
rect 5825 125 5835 181
rect 9035 125 9087 181
rect 5825 118 9087 125
rect 9041 77 9087 118
rect 9041 -164 9087 -123
rect 5825 -171 9087 -164
rect 5825 -227 5835 -171
rect 9035 -227 9087 -171
rect 9237 -368 9283 854
rect 9311 657 9321 713
rect 12521 657 12531 713
rect 9311 650 12531 657
rect 12755 696 12801 854
rect 13013 696 13059 854
rect 12755 650 12830 696
rect 12992 650 13059 696
rect 12517 409 12527 609
rect 12579 409 12589 609
rect 12755 368 12801 650
rect 13013 368 13059 650
rect 9311 361 12531 368
rect 9311 305 9321 361
rect 12521 305 12531 361
rect 12755 322 12831 368
rect 12995 322 13059 368
rect 9311 125 9321 181
rect 12521 125 12531 181
rect 9311 118 12531 125
rect 12755 164 12801 322
rect 13013 164 13059 322
rect 12755 118 12829 164
rect 12993 118 13059 164
rect 12517 -123 12527 77
rect 12579 -123 12589 77
rect 12755 -164 12801 118
rect 13013 -164 13059 118
rect 9311 -171 12531 -164
rect 9311 -227 9321 -171
rect 12521 -227 12531 -171
rect 12755 -210 12834 -164
rect 12990 -210 13059 -164
rect 12755 -368 12801 -210
rect 13013 -368 13059 -210
rect 1811 -414 13059 -368
rect 1811 -696 1857 -414
rect 2069 -696 2115 -414
rect 2265 -696 2343 -414
rect 5555 -696 5601 -414
rect 5751 -696 5829 -414
rect 9041 -696 9087 -414
rect 9237 -696 9315 -414
rect 12527 -696 12573 -414
rect 12755 -696 12801 -414
rect 13013 -696 13059 -414
rect 1811 -742 13059 -696
rect 13758 1182 13826 1228
rect 14004 1182 14062 1228
rect 13758 900 13804 1182
rect 14016 900 14062 1182
rect 13758 854 13828 900
rect 14004 854 14062 900
rect 13758 696 13804 854
rect 14016 696 14062 854
rect 13758 650 13824 696
rect 13994 650 14062 696
rect 13758 368 13804 650
rect 14016 368 14062 650
rect 13758 322 13826 368
rect 14003 322 14062 368
rect 13758 164 13804 322
rect 14016 164 14062 322
rect 13758 118 13822 164
rect 14001 118 14062 164
rect 13758 -164 13804 118
rect 14016 -164 14062 118
rect 13758 -210 13824 -164
rect 13998 -210 14062 -164
rect 13758 -368 13804 -210
rect 14016 -368 14062 -210
rect 14190 -368 14258 1918
rect 14286 1721 14296 1778
rect 15896 1721 15906 1778
rect 14286 1714 15906 1721
rect 16130 1760 16176 1918
rect 16388 1760 16434 1918
rect 16130 1714 16199 1760
rect 16374 1714 16434 1760
rect 15892 1473 15902 1673
rect 15954 1473 15964 1673
rect 16130 1432 16176 1714
rect 16388 1432 16434 1714
rect 14286 1425 15906 1432
rect 14286 1368 14296 1425
rect 15896 1368 15906 1425
rect 16130 1386 16200 1432
rect 16377 1386 16434 1432
rect 14286 1189 14296 1246
rect 15896 1189 15948 1246
rect 14286 1182 15948 1189
rect 15902 1140 15948 1182
rect 16130 1228 16176 1386
rect 16388 1228 16434 1386
rect 16130 1182 16194 1228
rect 16375 1182 16434 1228
rect 15902 900 15948 941
rect 14287 893 15948 900
rect 14287 836 14297 893
rect 15897 836 15948 893
rect 16130 900 16176 1182
rect 16388 900 16434 1182
rect 16130 854 16197 900
rect 16375 854 16434 900
rect 14286 657 14296 714
rect 15896 657 15948 714
rect 14286 650 15948 657
rect 15902 609 15948 650
rect 16130 696 16176 854
rect 16388 696 16434 854
rect 16130 650 16198 696
rect 16374 650 16434 696
rect 15902 368 15948 409
rect 14286 361 15948 368
rect 14286 304 14296 361
rect 15896 304 15948 361
rect 16130 368 16176 650
rect 16388 368 16434 650
rect 16130 322 16198 368
rect 16376 322 16434 368
rect 14286 125 14296 182
rect 15896 125 15906 182
rect 14286 118 15906 125
rect 16130 164 16176 322
rect 16388 164 16434 322
rect 16130 118 16195 164
rect 16370 118 16434 164
rect 15892 -123 15902 77
rect 15954 -123 15964 77
rect 16130 -164 16176 118
rect 16388 -164 16434 118
rect 14286 -171 15906 -164
rect 14286 -228 14296 -171
rect 15896 -228 15906 -171
rect 16130 -210 16200 -164
rect 16367 -210 16434 -164
rect 16130 -368 16176 -210
rect 16388 -368 16434 -210
rect 17478 -282 17678 -82
rect 13758 -414 16434 -368
rect 13758 -696 13804 -414
rect 14016 -696 14062 -414
rect 14190 -696 14291 -414
rect 15902 -696 15948 -414
rect 16130 -696 16176 -414
rect 16388 -696 16434 -414
rect 17478 -682 17678 -482
rect 13758 -742 16434 -696
rect 17478 -1082 17678 -882
rect 17478 -1482 17678 -1282
rect 14049 -1655 14095 -1654
rect 16725 -1655 16771 -1654
rect 13791 -1701 16771 -1655
rect 13791 -1965 13837 -1701
rect 14049 -1965 14095 -1701
rect 14429 -1965 14475 -1701
rect 16087 -1965 16133 -1701
rect 16467 -1965 16513 -1701
rect 16725 -1965 16771 -1701
rect 17478 -1882 17678 -1682
rect 13791 -2011 16771 -1965
rect 13791 -2241 13837 -2011
rect 14049 -2241 14095 -2011
rect 13791 -2287 13854 -2241
rect 14038 -2287 14095 -2241
rect 14471 -2271 14481 -2219
rect 16081 -2271 16091 -2219
rect 14471 -2287 16091 -2271
rect 16467 -2241 16513 -2011
rect 16725 -2241 16771 -2011
rect 16467 -2287 16530 -2241
rect 16710 -2287 16771 -2241
rect 17478 -2282 17678 -2082
rect 13791 -2611 13837 -2287
rect 14049 -2611 14095 -2287
rect 14413 -2579 14423 -2319
rect 14475 -2579 14485 -2319
rect 13791 -2657 13853 -2611
rect 14031 -2657 14095 -2611
rect 13791 -2887 13837 -2657
rect 14049 -2887 14095 -2657
rect 14471 -2627 16091 -2611
rect 14471 -2679 14481 -2627
rect 16081 -2679 16091 -2627
rect 13791 -2933 13854 -2887
rect 14032 -2933 14095 -2887
rect 14471 -2917 14481 -2865
rect 16081 -2917 16091 -2865
rect 14471 -2933 16091 -2917
rect 13791 -3257 13837 -2933
rect 14049 -3257 14095 -2933
rect 14413 -3225 14423 -2965
rect 14475 -3225 14485 -2965
rect 13791 -3303 13847 -3257
rect 14038 -3303 14095 -3257
rect 13791 -3533 13837 -3303
rect 14049 -3533 14095 -3303
rect 14471 -3325 14481 -3273
rect 16081 -3325 16091 -3273
rect 13791 -3579 13850 -3533
rect 14037 -3579 14095 -3533
rect 14471 -3563 14481 -3511
rect 16081 -3563 16091 -3511
rect 13791 -3903 13837 -3579
rect 14049 -3903 14095 -3579
rect 14413 -3871 14423 -3611
rect 14475 -3871 14485 -3611
rect 13791 -3949 13852 -3903
rect 14034 -3949 14095 -3903
rect 13791 -4179 13837 -3949
rect 14049 -4179 14095 -3949
rect 14471 -3919 16091 -3903
rect 14471 -3971 14481 -3919
rect 16081 -3971 16091 -3919
rect 13791 -4225 13847 -4179
rect 14038 -4225 14095 -4179
rect 14471 -4209 14481 -4157
rect 16081 -4209 16091 -4157
rect 14471 -4225 16091 -4209
rect 8939 -4389 9007 -4337
rect 13007 -4389 13017 -4337
rect 8939 -4405 13017 -4389
rect 8939 -4437 9011 -4405
rect 8939 -4637 8949 -4437
rect 9001 -4637 9011 -4437
rect 8939 -4669 9011 -4637
rect 8939 -4685 13017 -4669
rect 8939 -4737 9007 -4685
rect 13007 -4737 13017 -4685
rect 8997 -4903 9007 -4851
rect 13007 -4903 13017 -4851
rect 8997 -4919 13017 -4903
rect 8939 -5151 8949 -4951
rect 9001 -5151 9011 -4951
rect 8997 -5199 13017 -5183
rect 8997 -5251 9007 -5199
rect 13007 -5251 13017 -5199
rect 13045 -5399 13091 -4437
rect 13791 -4549 13837 -4225
rect 14049 -4549 14095 -4225
rect 14413 -4517 14423 -4257
rect 14475 -4517 14485 -4257
rect 16119 -4517 16165 -2319
rect 16467 -2611 16513 -2287
rect 16725 -2611 16771 -2287
rect 16467 -2657 16530 -2611
rect 16710 -2657 16771 -2611
rect 16467 -2887 16513 -2657
rect 16725 -2887 16771 -2657
rect 17478 -2682 17678 -2482
rect 16467 -2933 16529 -2887
rect 16708 -2933 16771 -2887
rect 16467 -3257 16513 -2933
rect 16725 -3257 16771 -2933
rect 16467 -3303 16529 -3257
rect 16712 -3303 16771 -3257
rect 16467 -3533 16513 -3303
rect 16725 -3533 16771 -3303
rect 16467 -3579 16528 -3533
rect 16714 -3579 16771 -3533
rect 16467 -3903 16513 -3579
rect 16725 -3903 16771 -3579
rect 16467 -3949 16527 -3903
rect 16712 -3949 16771 -3903
rect 16467 -4179 16513 -3949
rect 16725 -4179 16771 -3949
rect 16467 -4225 16530 -4179
rect 16710 -4225 16771 -4179
rect 16467 -4549 16513 -4225
rect 16725 -4549 16771 -4225
rect 13791 -4595 13850 -4549
rect 14037 -4595 14095 -4549
rect 13791 -4825 13837 -4595
rect 14049 -4825 14095 -4595
rect 14471 -4565 16091 -4549
rect 14471 -4617 14481 -4565
rect 16081 -4617 16091 -4565
rect 16467 -4595 16528 -4549
rect 16715 -4595 16771 -4549
rect 16467 -4825 16513 -4595
rect 16725 -4825 16771 -4595
rect 13791 -4871 16771 -4825
rect 13791 -5135 13837 -4871
rect 14049 -5135 14095 -4871
rect 14429 -5135 14475 -4871
rect 16087 -5135 16133 -4871
rect 16467 -5135 16513 -4871
rect 16725 -5135 16771 -4871
rect 13791 -5181 16771 -5135
rect 16467 -5182 16513 -5181
<< via1 >>
rect 2349 657 5549 713
rect 5555 409 5607 609
rect 2349 305 5549 361
rect 2349 125 5549 181
rect 5555 -123 5607 77
rect 2349 -227 5549 -171
rect 5835 657 9035 713
rect 5835 305 9035 361
rect 5835 125 9035 181
rect 5835 -227 9035 -171
rect 9321 657 12521 713
rect 12527 409 12579 609
rect 9321 305 12521 361
rect 9321 125 12521 181
rect 12527 -123 12579 77
rect 9321 -227 12521 -171
rect 14296 1721 15896 1778
rect 15902 1473 15954 1673
rect 14296 1368 15896 1425
rect 14296 1189 15896 1246
rect 14297 836 15897 893
rect 14296 657 15896 714
rect 14296 304 15896 361
rect 14296 125 15896 182
rect 15902 -123 15954 77
rect 14296 -228 15896 -171
rect 14481 -2271 16081 -2219
rect 14423 -2579 14475 -2319
rect 14481 -2679 16081 -2627
rect 14481 -2917 16081 -2865
rect 14423 -3225 14475 -2965
rect 14481 -3325 16081 -3273
rect 14481 -3563 16081 -3511
rect 14423 -3871 14475 -3611
rect 14481 -3971 16081 -3919
rect 14481 -4209 16081 -4157
rect 9007 -4389 13007 -4337
rect 8949 -4637 9001 -4437
rect 9007 -4737 13007 -4685
rect 9007 -4903 13007 -4851
rect 8949 -5151 9001 -4951
rect 9007 -5251 13007 -5199
rect 14423 -4517 14475 -4257
rect 14481 -4617 16081 -4565
<< metal2 >>
rect 13457 1781 16735 1791
rect 13614 1778 16578 1781
rect 13614 1721 14296 1778
rect 15896 1721 16578 1778
rect 13457 1711 16735 1721
rect 15902 1673 16974 1683
rect 15954 1473 16823 1673
rect 16964 1473 16974 1673
rect 15902 1463 16974 1473
rect 13457 1425 16735 1435
rect 13614 1368 14296 1425
rect 15896 1368 16578 1425
rect 13614 1365 16578 1368
rect 13457 1355 16735 1365
rect 13457 1249 16735 1259
rect 13614 1246 16578 1249
rect 13614 1189 14296 1246
rect 15896 1189 16578 1246
rect 13457 1179 16735 1189
rect 13457 893 16735 903
rect 5504 833 13457 836
rect 13614 836 14297 893
rect 15897 836 16578 893
rect 13614 833 16578 836
rect 5504 826 16735 833
rect 5661 766 12471 826
rect 12628 823 16735 826
rect 12628 766 13624 823
rect 5504 756 13624 766
rect 13457 727 13624 756
rect 2349 717 13377 727
rect 2349 713 13220 717
rect 5549 657 5835 713
rect 9035 657 9321 713
rect 12521 657 13220 713
rect 2349 647 13377 657
rect 13457 717 16735 727
rect 13614 714 16578 717
rect 13614 657 14296 714
rect 15896 657 16578 714
rect 13457 647 16735 657
rect 5553 609 5609 619
rect 5553 399 5609 409
rect 12525 609 12581 619
rect 12525 399 12581 409
rect 2349 361 13377 371
rect 5549 305 5835 361
rect 9035 305 9321 361
rect 12521 305 13220 361
rect 2349 301 13220 305
rect 2349 291 13377 301
rect 13457 361 16735 371
rect 13614 304 14296 361
rect 15896 304 16578 361
rect 13614 301 16578 304
rect 13457 291 16735 301
rect 2349 185 13377 195
rect 2349 181 13220 185
rect 5549 125 5835 181
rect 9035 125 9321 181
rect 12521 125 13220 181
rect 2349 115 13377 125
rect 13457 185 16735 195
rect 13614 182 16578 185
rect 13614 125 14296 182
rect 15896 125 16578 182
rect 13457 115 16735 125
rect 5553 77 5609 87
rect 5553 -133 5609 -123
rect 12525 77 12581 87
rect 12525 -133 12581 -123
rect 15902 77 16974 87
rect 15954 76 16974 77
rect 15954 -123 16822 76
rect 15902 -124 16822 -123
rect 16963 -124 16974 76
rect 15902 -133 16974 -124
rect 2349 -171 13377 -161
rect 5549 -227 5835 -171
rect 9035 -227 9321 -171
rect 12521 -227 13220 -171
rect 2349 -231 13220 -227
rect 2349 -241 13377 -231
rect 13457 -171 16735 -161
rect 13614 -228 14296 -171
rect 15896 -228 16577 -171
rect 13614 -231 16577 -228
rect 16734 -231 16735 -171
rect 13457 -241 16735 -231
rect 5504 -279 13614 -269
rect 5661 -339 12471 -279
rect 12628 -339 13457 -279
rect 5504 -349 13614 -339
rect 14183 -2209 14340 -2205
rect 14177 -2215 16081 -2209
rect 14177 -2275 14183 -2215
rect 14340 -2219 16081 -2215
rect 14340 -2271 14481 -2219
rect 14340 -2275 16081 -2271
rect 14177 -2281 16081 -2275
rect 14183 -2285 14340 -2281
rect 14421 -2319 14477 -2309
rect 14421 -2589 14477 -2579
rect 14183 -2617 14340 -2613
rect 14177 -2623 16081 -2617
rect 14177 -2683 14183 -2623
rect 14340 -2627 16081 -2623
rect 14340 -2679 14481 -2627
rect 14340 -2683 16081 -2679
rect 14177 -2689 16081 -2683
rect 14183 -2693 14340 -2689
rect 13447 -2742 14578 -2732
rect 13447 -2802 13457 -2742
rect 13614 -2802 14421 -2742
rect 13447 -2812 14578 -2802
rect 16221 -2855 16378 -2851
rect 14481 -2861 16385 -2855
rect 14481 -2865 16221 -2861
rect 16081 -2917 16221 -2865
rect 14481 -2921 16221 -2917
rect 16378 -2921 16385 -2861
rect 14481 -2927 16385 -2921
rect 16221 -2931 16378 -2927
rect 14421 -2965 14477 -2955
rect 14421 -3235 14477 -3225
rect 16221 -3263 16378 -3259
rect 14481 -3269 16385 -3263
rect 14481 -3273 16221 -3269
rect 16081 -3325 16221 -3273
rect 14481 -3329 16221 -3325
rect 16378 -3329 16385 -3269
rect 14481 -3335 16385 -3329
rect 16221 -3339 16378 -3335
rect 13210 -3388 14578 -3378
rect 13210 -3448 13220 -3388
rect 13377 -3448 14421 -3388
rect 13210 -3458 14578 -3448
rect 16221 -3501 16378 -3497
rect 14481 -3507 16385 -3501
rect 14481 -3511 16221 -3507
rect 16081 -3563 16221 -3511
rect 14481 -3567 16221 -3563
rect 16378 -3567 16385 -3507
rect 14481 -3573 16385 -3567
rect 16221 -3577 16378 -3573
rect 14421 -3611 14477 -3601
rect 14421 -3881 14477 -3871
rect 16221 -3909 16378 -3905
rect 14481 -3915 16385 -3909
rect 14481 -3919 16221 -3915
rect 16081 -3971 16221 -3919
rect 14481 -3975 16221 -3971
rect 16378 -3975 16385 -3915
rect 14481 -3981 16385 -3975
rect 16221 -3985 16378 -3981
rect 13210 -4034 14578 -4024
rect 13210 -4094 13220 -4034
rect 13377 -4094 14421 -4034
rect 13210 -4104 14578 -4094
rect 14183 -4147 14340 -4144
rect 14177 -4154 16081 -4147
rect 14177 -4214 14183 -4154
rect 14340 -4157 16081 -4154
rect 14340 -4209 14481 -4157
rect 14340 -4214 16081 -4209
rect 14177 -4219 16081 -4214
rect 14183 -4224 14340 -4219
rect 14421 -4257 14477 -4247
rect 8570 -4327 8727 -4323
rect 8560 -4333 13007 -4327
rect 8560 -4393 8570 -4333
rect 8727 -4337 13007 -4333
rect 8727 -4389 9007 -4337
rect 8727 -4393 13007 -4389
rect 8560 -4399 13007 -4393
rect 8570 -4403 8727 -4399
rect 8949 -4437 9001 -4427
rect 14421 -4527 14477 -4517
rect 14183 -4555 14340 -4551
rect 14183 -4561 16081 -4555
rect 14340 -4565 16081 -4561
rect 14340 -4617 14481 -4565
rect 14340 -4621 16081 -4617
rect 14183 -4627 16081 -4621
rect 14183 -4631 14340 -4627
rect 8949 -4647 9001 -4637
rect 8570 -4675 8727 -4671
rect 8560 -4681 13007 -4675
rect 8560 -4741 8570 -4681
rect 8727 -4685 13007 -4681
rect 8727 -4737 9007 -4685
rect 8727 -4741 13007 -4737
rect 8560 -4747 13007 -4741
rect 13447 -4680 14578 -4670
rect 13447 -4682 14421 -4680
rect 13447 -4742 13457 -4682
rect 13614 -4740 14421 -4682
rect 13614 -4742 14578 -4740
rect 8570 -4751 8727 -4747
rect 13447 -4750 14578 -4742
rect 8570 -4841 8727 -4837
rect 8560 -4847 13007 -4841
rect 8560 -4907 8570 -4847
rect 8727 -4851 13007 -4847
rect 8727 -4903 9007 -4851
rect 8727 -4907 13007 -4903
rect 8560 -4913 13007 -4907
rect 8570 -4917 8727 -4913
rect 8947 -4951 9003 -4941
rect 8947 -5161 9003 -5151
rect 8570 -5189 8727 -5185
rect 8560 -5195 13007 -5189
rect 8560 -5255 8570 -5195
rect 8727 -5199 13007 -5195
rect 8727 -5251 9007 -5199
rect 8727 -5255 13007 -5251
rect 8560 -5261 13007 -5255
rect 8570 -5265 8727 -5261
<< via2 >>
rect 13457 1721 13614 1781
rect 16578 1721 16735 1781
rect 16823 1473 16964 1673
rect 13457 1365 13614 1425
rect 16578 1365 16735 1425
rect 13457 1189 13614 1249
rect 16578 1189 16735 1249
rect 13457 833 13614 893
rect 16578 833 16735 893
rect 5504 766 5661 826
rect 12471 766 12628 826
rect 13220 657 13377 717
rect 13457 657 13614 717
rect 16578 657 16735 717
rect 5553 409 5555 609
rect 5555 409 5607 609
rect 5607 409 5609 609
rect 12525 409 12527 609
rect 12527 409 12579 609
rect 12579 409 12581 609
rect 13220 301 13377 361
rect 13457 301 13614 361
rect 16578 301 16735 361
rect 13220 125 13377 185
rect 13457 125 13614 185
rect 16578 125 16735 185
rect 5553 -123 5555 77
rect 5555 -123 5607 77
rect 5607 -123 5609 77
rect 12525 -123 12527 77
rect 12527 -123 12579 77
rect 12579 -123 12581 77
rect 16822 -124 16963 76
rect 13220 -231 13377 -171
rect 13457 -231 13614 -171
rect 16577 -231 16734 -171
rect 5504 -339 5661 -279
rect 12471 -339 12628 -279
rect 13457 -339 13614 -279
rect 14183 -2275 14340 -2215
rect 14421 -2579 14423 -2319
rect 14423 -2579 14475 -2319
rect 14475 -2579 14477 -2319
rect 14183 -2683 14340 -2623
rect 13457 -2802 13614 -2742
rect 14421 -2802 14578 -2742
rect 16221 -2921 16378 -2861
rect 14421 -3225 14423 -2965
rect 14423 -3225 14475 -2965
rect 14475 -3225 14477 -2965
rect 16221 -3329 16378 -3269
rect 13220 -3448 13377 -3388
rect 14421 -3448 14578 -3388
rect 16221 -3567 16378 -3507
rect 14421 -3871 14423 -3611
rect 14423 -3871 14475 -3611
rect 14475 -3871 14477 -3611
rect 16221 -3975 16378 -3915
rect 13220 -4094 13377 -4034
rect 14421 -4094 14578 -4034
rect 14183 -4214 14340 -4154
rect 8570 -4393 8727 -4333
rect 14421 -4517 14423 -4257
rect 14423 -4517 14475 -4257
rect 14475 -4517 14477 -4257
rect 14183 -4621 14340 -4561
rect 8570 -4741 8727 -4681
rect 13457 -4742 13614 -4682
rect 14421 -4740 14578 -4680
rect 8570 -4907 8727 -4847
rect 8947 -5151 8949 -4951
rect 8949 -5151 9001 -4951
rect 9001 -5151 9003 -4951
rect 8570 -5255 8727 -5195
<< metal3 >>
rect 13447 1781 13624 1792
rect 13447 1721 13457 1781
rect 13614 1721 13624 1781
rect 13447 1425 13624 1721
rect 13447 1365 13457 1425
rect 13614 1365 13624 1425
rect 13447 1249 13624 1365
rect 13447 1189 13457 1249
rect 13614 1189 13624 1249
rect 13447 893 13624 1189
rect 13447 833 13457 893
rect 13614 833 13624 893
rect 5494 826 5671 831
rect 5494 766 5504 826
rect 5661 766 5671 826
rect 5494 761 5671 766
rect 12461 826 12638 831
rect 12461 766 12471 826
rect 12628 766 12638 826
rect 12461 761 12638 766
rect 5543 609 5619 761
rect 5543 409 5553 609
rect 5609 409 5619 609
rect 5543 77 5619 409
rect 5543 -123 5553 77
rect 5609 -123 5619 77
rect 5543 -274 5619 -123
rect 12515 609 12591 761
rect 12515 409 12525 609
rect 12581 409 12591 609
rect 12515 77 12591 409
rect 12515 -123 12525 77
rect 12581 -123 12591 77
rect 12515 -274 12591 -123
rect 13210 717 13387 728
rect 13210 657 13220 717
rect 13377 657 13387 717
rect 13210 361 13387 657
rect 13210 301 13220 361
rect 13377 301 13387 361
rect 13210 185 13387 301
rect 13210 125 13220 185
rect 13377 125 13387 185
rect 13210 -171 13387 125
rect 13210 -231 13220 -171
rect 13377 -231 13387 -171
rect 13210 -236 13387 -231
rect 13447 717 13624 833
rect 13447 657 13457 717
rect 13614 657 13624 717
rect 13447 361 13624 657
rect 13447 301 13457 361
rect 13614 301 13624 361
rect 13447 185 13624 301
rect 13447 125 13457 185
rect 13614 125 13624 185
rect 13447 -171 13624 125
rect 13447 -231 13457 -171
rect 13614 -231 13624 -171
rect 5494 -279 5671 -274
rect 5494 -339 5504 -279
rect 5661 -339 5671 -279
rect 5494 -344 5671 -339
rect 12461 -279 12638 -274
rect 12461 -339 12471 -279
rect 12628 -339 12638 -279
rect 12461 -344 12638 -339
rect 13447 -279 13624 -231
rect 16567 1781 16745 1791
rect 16567 1721 16578 1781
rect 16735 1721 16745 1781
rect 16567 1425 16745 1721
rect 16567 1365 16578 1425
rect 16735 1365 16745 1425
rect 16567 1249 16745 1365
rect 16567 1189 16578 1249
rect 16735 1189 16745 1249
rect 16567 893 16745 1189
rect 16567 833 16578 893
rect 16735 833 16745 893
rect 16567 717 16745 833
rect 16567 657 16578 717
rect 16735 657 16745 717
rect 16567 361 16745 657
rect 16567 301 16578 361
rect 16735 301 16745 361
rect 16567 185 16745 301
rect 16567 125 16578 185
rect 16735 125 16745 185
rect 16567 -171 16745 125
rect 16567 -231 16577 -171
rect 16734 -231 16745 -171
rect 16567 -241 16745 -231
rect 16805 1673 16974 1683
rect 16805 1473 16823 1673
rect 16964 1473 16974 1673
rect 16805 76 16974 1473
rect 16805 -124 16822 76
rect 16963 -124 16974 76
rect 16805 -236 16974 -124
rect 13447 -339 13457 -279
rect 13614 -339 13624 -279
rect 13447 -375 13624 -339
rect 13210 -3388 13387 -2207
rect 13210 -3448 13220 -3388
rect 13377 -3448 13387 -3388
rect 13210 -4034 13387 -3448
rect 13210 -4094 13220 -4034
rect 13377 -4094 13387 -4034
rect 13210 -4104 13387 -4094
rect 13447 -2742 13624 -1733
rect 13447 -2802 13457 -2742
rect 13614 -2802 13624 -2742
rect 8560 -4333 8737 -4241
rect 8560 -4393 8570 -4333
rect 8727 -4393 8737 -4333
rect 8560 -4681 8737 -4393
rect 8560 -4741 8570 -4681
rect 8727 -4741 8737 -4681
rect 8560 -4847 8737 -4741
rect 13447 -4682 13624 -2802
rect 13447 -4742 13457 -4682
rect 13614 -4742 13624 -4682
rect 13447 -4750 13624 -4742
rect 14173 -2215 14350 -2210
rect 14173 -2275 14183 -2215
rect 14340 -2275 14350 -2215
rect 14173 -2623 14350 -2275
rect 14173 -2683 14183 -2623
rect 14340 -2683 14350 -2623
rect 14173 -4154 14350 -2683
rect 14411 -2319 14487 -2314
rect 14411 -2579 14421 -2319
rect 14477 -2579 14487 -2319
rect 14411 -2737 14487 -2579
rect 14411 -2742 14588 -2737
rect 14411 -2802 14421 -2742
rect 14578 -2802 14588 -2742
rect 14411 -2807 14588 -2802
rect 16211 -2861 16388 -2856
rect 16211 -2921 16221 -2861
rect 16378 -2921 16388 -2861
rect 14411 -2965 14487 -2960
rect 14411 -3225 14421 -2965
rect 14477 -3225 14487 -2965
rect 14411 -3383 14487 -3225
rect 16211 -3269 16388 -2921
rect 16211 -3329 16221 -3269
rect 16378 -3329 16388 -3269
rect 14411 -3388 14588 -3383
rect 14411 -3448 14421 -3388
rect 14578 -3448 14588 -3388
rect 14411 -3453 14588 -3448
rect 16211 -3507 16388 -3329
rect 16211 -3567 16221 -3507
rect 16378 -3567 16388 -3507
rect 14411 -3611 14487 -3606
rect 14411 -3871 14421 -3611
rect 14477 -3871 14487 -3611
rect 14411 -4029 14487 -3871
rect 16211 -3915 16388 -3567
rect 16211 -3975 16221 -3915
rect 16378 -3975 16388 -3915
rect 14411 -4034 14588 -4029
rect 14411 -4094 14421 -4034
rect 14578 -4094 14588 -4034
rect 14411 -4099 14588 -4094
rect 14173 -4214 14183 -4154
rect 14340 -4214 14350 -4154
rect 14173 -4561 14350 -4214
rect 14173 -4621 14183 -4561
rect 14340 -4621 14350 -4561
rect 8560 -4907 8570 -4847
rect 8727 -4907 8737 -4847
rect 8560 -5195 8737 -4907
rect 8560 -5255 8570 -5195
rect 8727 -5255 8737 -5195
rect 8560 -5261 8737 -5255
rect 8937 -4951 9013 -4946
rect 8937 -5151 8947 -4951
rect 9003 -5151 9013 -4951
rect 8937 -5610 9013 -5151
rect 14173 -5452 14350 -4621
rect 14411 -4257 14487 -4252
rect 14411 -4517 14421 -4257
rect 14477 -4517 14487 -4257
rect 14411 -4675 14487 -4517
rect 14411 -4680 14588 -4675
rect 14411 -4740 14421 -4680
rect 14578 -4740 14588 -4680
rect 14411 -4745 14588 -4740
rect 16211 -5390 16388 -3975
use trans_gate  x1
timestamp 1712344797
transform 1 0 3949 0 1 -2291
box 0 -2052 3413 715
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[0]
timestamp 1712597941
transform 1 0 15281 0 1 -2449
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM1[1]
timestamp 1712597941
transform 1 0 15281 0 1 -4387
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[0]
timestamp 1712597941
transform 1 0 15281 0 1 -3095
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_6975WM  XM2[1]
timestamp 1712597941
transform 1 0 15281 0 1 -3741
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[0]
timestamp 1712343889
transform 1 0 15096 0 1 1041
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM3[1]
timestamp 1712343889
transform 1 0 15096 0 1 509
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM4[0]
timestamp 1712669456
transform 1 0 7435 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1712671997
transform 1 0 7435 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[0]
timestamp 1712343889
transform 1 0 15096 0 1 1573
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM5[1]
timestamp 1712343889
transform 1 0 15096 0 1 -23
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[0]
timestamp 1712669456
transform 1 0 3949 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1712671997
transform 1 0 3949 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_CDT3CS  XM6[2]
timestamp 1712669456
transform 1 0 10921 0 1 509
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1712671997
transform 1 0 10921 0 1 -23
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1712343889
transform 1 0 11214 0 1 -1896
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_697RXD  XM8
timestamp 1712343889
transform 1 0 11184 0 1 -2752
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1712343889
transform 1 0 12907 0 1 -1704
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1712343889
transform 1 0 12907 0 1 -2883
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1712343889
transform 1 0 11007 0 1 -4537
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1712343889
transform 1 0 11007 0 1 -5051
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1712343889
transform 1 0 9394 0 1 -2732
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1712343889
transform 1 0 9394 0 1 -3459
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1712343889
transform 1 0 12397 0 1 2117
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1712343889
transform 1 0 11109 0 1 2136
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1712343889
transform 1 0 10714 0 1 -3505
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1712343889
transform 1 0 8258 0 1 -1892
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1712343889
transform 1 0 8260 0 1 -2732
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[0]
timestamp 1712671997
transform 1 0 13910 0 1 2105
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[1]
timestamp 1712671997
transform 1 0 13910 0 1 1573
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[2]
timestamp 1712671997
transform 1 0 13910 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[3]
timestamp 1712671997
transform 1 0 13910 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712671997
transform 1 0 13910 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712671997
transform 1 0 13910 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712671997
transform 1 0 16282 0 1 2105
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712671997
transform 1 0 16282 0 1 1573
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712671997
transform 1 0 16282 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712671997
transform 1 0 16282 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712671997
transform 1 0 16282 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712671997
transform 1 0 16282 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712671997
transform 1 0 1963 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712671997
transform 1 0 1963 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712671997
transform 1 0 1963 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712671997
transform 1 0 1963 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[16]
timestamp 1712671997
transform 1 0 12907 0 1 1041
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[17]
timestamp 1712671997
transform 1 0 12907 0 1 509
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[18]
timestamp 1712671997
transform 1 0 12907 0 1 -23
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[19]
timestamp 1712671997
transform 1 0 12907 0 1 -555
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[0]
timestamp 1712343889
transform 1 0 15096 0 1 2105
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD8[1]
timestamp 1712343889
transform 1 0 15096 0 1 -555
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712671997
transform 1 0 3949 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712671997
transform 1 0 7435 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712671997
transform 1 0 10921 0 1 1041
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712671997
transform 1 0 3949 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712671997
transform 1 0 7435 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712671997
transform 1 0 10921 0 1 -555
box -1796 -319 1796 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712600458
transform 1 0 13943 0 1 -1833
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712600458
transform 1 0 13943 0 1 -5003
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712600458
transform 1 0 16619 0 1 -1833
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712600458
transform 1 0 16619 0 1 -5003
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712599722
transform 1 0 15281 0 1 -1833
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712599722
transform 1 0 15281 0 1 -5003
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712597941
transform 1 0 13943 0 1 -2449
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712597941
transform 1 0 13943 0 1 -3095
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712597941
transform 1 0 13943 0 1 -3741
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712597941
transform 1 0 13943 0 1 -4387
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[4]
timestamp 1712597941
transform 1 0 16619 0 1 -2449
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[5]
timestamp 1712597941
transform 1 0 16619 0 1 -3095
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[6]
timestamp 1712597941
transform 1 0 16619 0 1 -3741
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[7]
timestamp 1712597941
transform 1 0 16619 0 1 -4387
box -328 -388 328 388
<< labels >>
flabel metal1 17478 -1882 17678 -1682 0 FreeSans 256 180 0 0 vref
port 2 nsew
flabel metal1 17478 -1482 17678 -1282 0 FreeSans 256 180 0 0 vin
port 3 nsew
flabel metal1 17478 -1082 17678 -882 0 FreeSans 256 180 0 0 ena
port 4 nsew
flabel metal1 17478 -682 17678 -482 0 FreeSans 256 180 0 0 ibias
port 5 nsew
flabel metal1 17478 -282 17678 -82 0 FreeSans 256 180 0 0 vss
port 6 nsew
flabel metal1 17478 -2282 17678 -2082 0 FreeSans 256 180 0 0 out
port 1 nsew
flabel metal1 17478 -2682 17678 -2482 0 FreeSans 256 180 0 0 dvdd
port 0 nsew
<< end >>

* NGSPICE file created from sky130_vbl_ip__overvoltage.ext - technology: sky130A

.subckt sky130_vbl_ip__overvoltage vtrip[3] vtrip[2] ovout vtrip[0] vbg ibias ena
+ vtrip[1] dvss dvdd avdd avss
X0 dvss.t67 dvss.t65 dvss.t66 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X1 multiplexer_0.trans_gate_m_31.out.t0 multiplexer_0.vtrip_1.t0 multiplexer_0.trans_gate_m_29.in.t3 avss.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X2 avss.t98 multiplexer_0.vtrip_1_b.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X3 a_n15874_n447# a_n12654_n447# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X4 a_n12118_12027# a_n8898_11649# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X5 dvss.t64 dvss.t62 dvss.t63 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X6 avss.t190 avss.t191 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X7 avss.t133 avss.t134 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X8 comp_hyst_0.net3.t0 comp_hyst_0.net4 dvdd.t118 dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X9 avss.t91 avss.t92 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X10 avss.t202 avss.t203 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X11 avss.t240 level_shifter_3.in_b.t2 multiplexer_0.vtrip_3.t0 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X12 a_n8362_4845# multiplexer_0.in_0110.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X13 a_n15874_8625# a_n12654_9003# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X14 avss.t19 multiplexer_0.vtrip_2.t1 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X15 a_n12118_9759# a_n8898_9381# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X16 multiplexer_0.in_1100.t3 multiplexer_0.in_1101.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X17 dvss.t61 dvss.t59 dvss.t60 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X18 a_n15874_6357# a_n12654_5979# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X19 level_shifter_0.in_b.t0 vtrip[0].t0 dvdd.t93 dvdd.t92 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X20 dvdd.t91 dvdd.t89 dvdd.t90 dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X21 multiplexer_0.trans_gate_m_37.out.t2 multiplexer_0.vtrip_2.t2 multiplexer_0.trans_gate_m_32.in.t1 avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X22 multiplexer_0.trans_gate_m_21.in.t1 multiplexer_0.vtrip_0.t0 multiplexer_0.in_1011.t2 avss.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X23 avss.t169 vtrip[1].t0 multiplexer_0.vtrip_1_b.t0 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X24 dvss.t4 comp_hyst_0.net5 comp_hyst_0.net1 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X25 avss.t159 avss.t160 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X26 multiplexer_0.trans_gate_m_29.in.t4 multiplexer_0.vtrip_0.t1 multiplexer_0.in_0010.t3 avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X27 avss.t95 multiplexer_0.vtrip_0_b.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X28 a_n12118_2955# a_n8898_3333# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X29 avss.t83 avss.t84 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X30 avss.t183 avss.t184 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X31 voltage_divider_0.51 multiplexer_0.in_0000.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X32 avss.t60 avss.t61 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X33 comp_hyst_0.net1.t1 comp_hyst_0.vin comp_hyst_0.net3.t0 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X34 a_n15874_13161# a_n12654_13539# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X35 multiplexer_0.trans_gate_m_23.in.t3 multiplexer_0.vtrip_0_b.t3 multiplexer_0.in_1001.t2 avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X36 a_n8362_13161# a_n5142_12783# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X37 avss.t172 avss.t173 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X38 avss.t157 avss.t158 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X39 a_n12118_7491# a_n8898_7113# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X40 multiplexer_0.trans_gate_m_32.in.t2 multiplexer_0.vtrip_1.t1 multiplexer_0.trans_gate_m_23.in.t4 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X41 multiplexer_0.vtrip_2.t0 multiplexer_0.vtrip_2_b.t2 avdd.t6 avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X42 avss.t89 avss.t90 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X43 dvdd.t88 dvdd.t86 dvdd.t87 dvdd.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X44 a_n15874_3333# a_n12654_3711# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X45 a_n8898_n447# a_n5142_n825# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X46 comp_hyst_0.net1.t2 vbg.t0 comp_hyst_0.net4 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X47 avss.t67 avss.t68 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X48 avss.t154 avss.t155 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X49 avss.t222 level_shifter_0.in_b.t2 level_shifter_0.out avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X50 a_n12118_10515# a_n8898_10893# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X51 comp_hyst_0.net4 comp_hyst_0.net3.t0 dvdd.t105 dvdd.t44 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X52 a_n8362_8625# multiplexer_0.in_0000.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X53 multiplexer_0.in_0100.t3 a_n5142_5979# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X54 dvdd.t85 dvdd.t83 dvdd.t84 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X55 a_n15874_10893# a_n12654_11271# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X56 comp_hyst_0.net1.t0 comp_hyst_0.vin comp_hyst_0.net3.t0 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X57 multiplexer_0.trans_gate_m_27.in.t1 multiplexer_0.vtrip_0.t2 multiplexer_0.in_0101.t2 avss.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X58 avss.t111 avss.t112 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X59 comp_hyst_0.net1.t3 vbg.t1 comp_hyst_0.net4 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X60 avss.t151 avss.t152 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X61 a_n8362_10137# a_n5142_9759# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X62 a_n12118_6735# a_n8898_7113# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X63 multiplexer_0.trans_gate_m_28.in.t4 multiplexer_0.vtrip_1_b.t3 multiplexer_0.trans_gate_m_27.in.t5 avss.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X64 avss.t224 ena.t0 a_n5142_n1959.t0 avss.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=3
X65 dvdd.t82 dvdd.t80 dvdd.t81 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X66 a_n12118_4467# a_n8898_4089# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X67 avss.t109 avss.t110 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X68 dvss.t58 dvss.t56 dvss.t57 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X69 a_n15874_1065# a_n12654_1065# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X70 multiplexer_0.vtrip_3.t1 multiplexer_0.vtrip_3_b.t2 avdd.t27 avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X71 vin.t3 multiplexer_0.vtrip_3_b.t3 multiplexer_0.trans_gate_m_33.in.t2 avss.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X72 avss.t185 multiplexer_0.vtrip_1_b.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X73 avss.t230 avss.t231 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X74 a_n8362_13917# a_n5142_14295# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X75 dvdd.t79 dvdd.t77 dvdd.t78 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X76 multiplexer_0.trans_gate_m_33.in.t3 multiplexer_0.vtrip_2.t3 multiplexer_0.trans_gate_m_31.out.t1 avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X77 avss.t126 avss.t127 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X78 a_n12118_10515# a_n8898_10137# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X79 avss.t179 avss.t180 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X80 a_n8362_13917# a_n5142_13539# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X81 multiplexer_0.in_1010.t1 multiplexer_0.in_1001.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X82 a_n15874_n447# a_n12654_n69# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X83 a_n15874_4845# a_n12654_4467# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X84 avss.t181 avss.t182 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X85 dvss.t13 comp_hyst_0.ena_b comp_hyst_0.net5.t2 dvss.t12 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X86 a_n12118_14295# a_n8898_14673# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X87 level_shifter_2.in_b.t0 vtrip[2].t0 dvdd.t110 dvdd.t109 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X88 dvdd.t76 dvdd.t74 dvdd.t75 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X89 a_n12654_1821# a_n8898_1821# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X90 a_n15874_14673# a_n12654_15051# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X91 avss.t124 avss.t125 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X92 multiplexer_0.trans_gate_m_18.in.t1 multiplexer_0.vtrip_0.t3 multiplexer_0.in_1100.t1 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X93 avss.t7 level_shifter_2.in_b.t2 level_shifter_2.out avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X94 avss.t30 avss.t31 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X95 multiplexer_0.trans_gate_m_32.in.t4 multiplexer_0.vtrip_1_b.t5 multiplexer_0.trans_gate_m_21.in.t4 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X96 comp_hyst_0.net3.t2 comp_hyst_0.net3.t0 dvdd.t104 dvdd.t26 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X97 avss.t54 avss.t55 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X98 dvss.t22 vtrip[2].t1 level_shifter_2.in_b.t1 dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X99 a_n12118_8247# a_n8898_7869# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X100 multiplexer_0.trans_gate_m_19.in.t2 multiplexer_0.vtrip_0_b.t4 multiplexer_0.in_1110.t1 avss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X101 dvss.t75 comp_hyst_0.net2 comp_hyst_0.net2 dvss.t74 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X102 a_n15874_n1959# a_n12654_n1959# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X103 a_n8898_1065# a_n5142_687# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X104 multiplexer_0.vtrip_0_b.t0 level_shifter_0.out avdd.t22 avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X105 multiplexer_0.trans_gate_m_29.in.t0 multiplexer_0.vtrip_0_b.t5 multiplexer_0.in_0011.t2 avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X106 avss.t28 avss.t29 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X107 multiplexer_0.trans_gate_m_33.in.t2 multiplexer_0.vtrip_2.t4 multiplexer_0.trans_gate_m_28.in.t1 avss.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X108 avss.t98 multiplexer_0.vtrip_1.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X109 dvdd.t73 dvdd.t71 dvdd.t72 dvdd.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X110 a_n8898_n1581# a_n5142_n1581# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X111 a_n15874_1821# a_n12654_2199# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X112 a_n12654_n69# a_n8898_n69# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X113 a_n12118_11271# a_n8898_11649# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X114 avss.t42 avss.t43 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X115 a_n8362_4845# multiplexer_0.in_0111.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X116 a_n15874_11649# a_n12654_12027# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X117 a_n15874_8625# a_n12654_8247# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X118 avss.t57 avss.t58 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X119 multiplexer_0.trans_gate_m_19.in.t1 multiplexer_0.vtrip_0.t4 multiplexer_0.in_1111.t0 avss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X120 avss.t177 avss.t178 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X121 a_n15874_5601# a_n12654_5979# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X122 avss.t95 multiplexer_0.vtrip_0.t5 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X123 multiplexer_0.trans_gate_m_28.in.t1 multiplexer_0.vtrip_1.t3 multiplexer_0.trans_gate_m_25.in.t4 avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X124 comp_hyst_0.net4 comp_hyst_0.net3.t0 dvdd.t103 dvdd.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X125 avss.t105 avss.t106 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X126 avss.t40 avss.t41 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X127 multiplexer_0.trans_gate_m_37.in.t2 multiplexer_0.vtrip_1.t4 multiplexer_0.trans_gate_m_19.in.t4 avss.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X128 a_n12118_5223# a_n8898_5601# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X129 a_n8898_n1203# a_n5142_n1581# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X130 a_n12118_2955# a_n8898_2577# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X131 avss.t248 avss.t249 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X132 multiplexer_0.trans_gate_m_25.in.t3 multiplexer_0.vtrip_0_b.t6 multiplexer_0.in_0111.t2 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X133 dvdd.t70 dvdd.t68 dvdd.t69 dvdd.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X134 avss.t228 avss.t229 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X135 comp_hyst_0.net4 ena.t1 dvdd.t120 dvdd.t119 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X136 avss.t26 avss.t27 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X137 a_n8362_12405# a_n5142_12783# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X138 multiplexer_0.trans_gate_m_23.in.t2 multiplexer_0.vtrip_0_b.t7 multiplexer_0.in_1000.t2 avss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X139 multiplexer_0.trans_gate_m_37.out.t1 multiplexer_0.vtrip_2_b.t3 multiplexer_0.trans_gate_m_37.in.t0 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X140 avss.t100 ena.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X141 dvdd.t67 dvdd.t65 dvdd.t66 dvdd.t44 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X142 multiplexer_0.in_1110.t3 multiplexer_0.in_1101.t2 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X143 dvdd.t64 dvdd.t62 dvdd.t63 dvdd.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X144 multiplexer_0.vtrip_3_b.t0 multiplexer_0.vtrip_3.t2 avdd.t17 avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X145 comp_hyst_0.net2 comp_hyst_0.net4 dvdd.t117 dvdd.t116 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X146 vin.t1 multiplexer_0.vtrip_3.t3 multiplexer_0.trans_gate_m_37.out.t4 avss.t227 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X147 avss.t65 avss.t66 avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X148 multiplexer_0.trans_gate_m_27.in.t0 multiplexer_0.vtrip_0.t6 multiplexer_0.in_0100.t1 avdd.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X149 avss.t255 avss.t256 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X150 avss.t81 avss.t82 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X151 avss.t46 avss.t47 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X152 multiplexer_0.trans_gate_m_31.in.t1 multiplexer_0.vtrip_0.t7 multiplexer_0.in_0000.t1 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X153 a_n8362_8625# multiplexer_0.in_0001.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X154 avss.t44 avss.t45 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X155 multiplexer_0.in_0101.t1 a_n5142_5979# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X156 multiplexer_0.trans_gate_m_37.in.t3 multiplexer_0.vtrip_1.t5 multiplexer_0.trans_gate_m_18.in.t4 avdd.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X157 a_n12654_n825# a_n8898_n825# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X158 avss.t101 avss.t102 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X159 a_n15874_9381# a_n12654_9759# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X160 a_n15874_10893# a_n12654_10515# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X161 avss.t170 avss.t171 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X162 a_n8362_12405# a_n5142_12027# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X163 dvss.t10 vbg.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X164 a_n12118_6735# a_n8898_6357# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X165 avss.t121 avss.t122 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X166 a_n15874_3333# a_n12654_2955# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X167 avss.t87 avss.t88 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X168 avss.t17 avss.t18 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X169 a_n12118_12783# a_n8898_13161# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X170 multiplexer_0.trans_gate_m_18.in.t2 multiplexer_0.vtrip_0_b.t8 multiplexer_0.in_1101.t0 avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X171 dvss.t69 comp_hyst_0.ena_b.t0 comp_hyst_0.net2 dvss.t68 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X172 dvdd.t61 dvdd.t59 dvdd.t60 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X173 multiplexer_0.trans_gate_m_31.out.t4 multiplexer_0.vtrip_1.t6 multiplexer_0.trans_gate_m_31.in.t4 avdd.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X174 a_n15874_7113# a_n12654_7491# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X175 comp_hyst_0.ena_b ena.t3 dvdd.t107 dvdd.t106 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X176 a_n15874_10137# a_n12654_10515# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X177 avss.t9 avss.t10 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X178 multiplexer_0.trans_gate_m_37.out.t0 multiplexer_0.vtrip_2_b.t4 multiplexer_0.trans_gate_m_32.in.t0 avss.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X179 level_shifter_1.out multiplexer_0.vtrip_1_b.t6 avdd.t37 avdd.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X180 avss.t119 avss.t120 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X181 multiplexer_0.trans_gate_m_29.in.t1 multiplexer_0.vtrip_0_b.t9 multiplexer_0.in_0010.t1 avss.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X182 dvdd.t58 dvdd.t56 dvdd.t57 dvdd.t26 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X183 a_n12118_3711# a_n8898_4089# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X184 avss.t129 multiplexer_0.vtrip_3_b.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X185 avss.t85 avss.t86 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X186 avss.t210 avss.t211 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X187 avss.t72 vtrip[3].t0 multiplexer_0.vtrip_3_b.t1 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X188 a_n15874_309# a_n12654_687# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X189 voltage_divider_0.51 a_n5142_9759# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X190 a_n15874_14673# a_n12654_14295# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X191 dvdd.t55 dvdd.t53 dvdd.t54 dvdd.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X192 dvss.t15 ena.t4 comp_hyst_0.ena_b dvss.t14 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X193 multiplexer_0.trans_gate_m_23.in.t1 multiplexer_0.vtrip_0.t8 multiplexer_0.in_1001.t1 avss.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X194 comp_hyst_0.net5 ena.t5 ibias.t1 dvss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
X195 a_n12118_9759# a_n8898_10137# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X196 avss.t141 avss.t142 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X197 a_n8362_13161# a_n5142_13539# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X198 multiplexer_0.trans_gate_m_32.in.t0 multiplexer_0.vtrip_1_b.t7 multiplexer_0.trans_gate_m_23.in.t5 avss.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X199 multiplexer_0.in_1010.t0 multiplexer_0.in_1011.t1 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X200 a_n15874_7113# a_n12654_6735# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X201 a_n12118_7491# a_n8898_7869# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X202 a_n15874_4089# a_n12654_4467# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X203 avss.t139 avss.t140 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X204 dvss.t11 ena.t6 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X205 a_n12118_14295# a_n8898_13917# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X206 level_shifter_1.in_b.t0 vtrip[1].t1 dvdd.t112 dvdd.t111 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X207 dvdd.t52 dvdd.t50 dvdd.t51 dvdd.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X208 avss.t117 avss.t118 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X209 multiplexer_0.trans_gate_m_21.in.t0 multiplexer_0.vtrip_0.t9 multiplexer_0.in_1010.t2 avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X210 dvdd.t49 dvdd.t47 dvdd.t48 dvdd.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X211 multiplexer_0.trans_gate_m_28.in.t2 multiplexer_0.vtrip_1.t7 multiplexer_0.trans_gate_m_27.in.t4 avdd.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X212 a_n12118_13539# a_n8898_13917# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X213 a_n12654_1443# a_n8898_1443# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X214 a_n8362_7113# multiplexer_0.in_0010.t2 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X215 avss.t63 avss.t64 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X216 avss.t69 level_shifter_1.in_b.t2 level_shifter_1.out avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X217 a_n15874_309# a_n12654_309# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X218 a_n8898_n69# a_n5142_n69# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X219 avss.t103 avss.t104 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X220 a_n12654_687# a_n8898_687# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X221 a_n15874_11649# a_n12654_11271# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X222 dvdd.t46 dvdd.t43 dvdd.t45 dvdd.t44 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X223 dvss.t1 vtrip[3].t1 level_shifter_3.in_b.t0 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X224 dvdd.t42 dvdd.t40 dvdd.t41 dvdd.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X225 a_n8362_10893# a_n5142_11271# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X226 avss.t79 avss.t80 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X227 avss.t220 avss.t221 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X228 multiplexer_0.trans_gate_m_18.in.t0 multiplexer_0.vtrip_0.t10 multiplexer_0.in_1101.t1 avss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X229 avss.t253 avss.t254 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X230 dvss.t7 vtrip[1].t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X231 avss.t38 avss.t39 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X232 dvdd.t39 dvdd.t36 dvdd.t38 dvdd.t37 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X233 a_n15874_1821# a_n12654_1821# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X234 comp_hyst_0.net4 comp_hyst_0.net3.t0 dvdd.t102 dvdd.t44 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X235 multiplexer_0.trans_gate_m_31.in.t2 multiplexer_0.vtrip_0_b.t10 multiplexer_0.in_0001.t3 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X236 avss.t36 avss.t37 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X237 multiplexer_0.trans_gate_m_25.in.t2 multiplexer_0.vtrip_0_b.t11 multiplexer_0.in_0110.t1 avss.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X238 avss.t245 avss.t246 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X239 multiplexer_0.trans_gate_m_33.in.t0 multiplexer_0.vtrip_2_b.t5 multiplexer_0.trans_gate_m_31.out.t0 avss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X240 multiplexer_0.trans_gate_m_37.in.t4 multiplexer_0.vtrip_1_b.t8 multiplexer_0.trans_gate_m_19.in.t5 avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X241 avss.t243 avss.t244 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X242 a_n8362_7113# multiplexer_0.in_0011.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X243 a_n12654_n1581# a_n8898_n1581# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X244 multiplexer_0.in_1000.t0 multiplexer_0.in_0111.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X245 a_n15874_7869# a_n12654_8247# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X246 dvss.t9 vtrip[1].t3 level_shifter_1.in_b.t1 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X247 a_n12654_309# a_n8898_309# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X248 comp_hyst_0.net4 comp_hyst_0.net4 dvdd.t115 dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X249 avss.t25 vtrip[0].t1 multiplexer_0.vtrip_0_b.t1 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X250 avss.t145 avss.t146 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X251 avss.t34 avss.t35 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X252 a_n12118_5223# a_n8898_4845# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X253 a_n12118_2199# a_n8898_2577# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X254 level_shifter_3.in_b.t1 vtrip[3].t2 dvdd.t97 dvdd.t96 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X255 avss.t217 avss.t218 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X256 dvdd.t35 dvdd.t33 dvdd.t34 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X257 multiplexer_0.trans_gate_m_31.out.t3 multiplexer_0.vtrip_1_b.t9 multiplexer_0.trans_gate_m_29.in.t2 avdd.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X258 avss.t131 multiplexer_0.vtrip_0.t11 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X259 a_n8898_15051# avdd.t19 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X260 avss.t241 avss.t242 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X261 avss.t215 avss.t216 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X262 avss.t14 avss.t15 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X263 avss.t115 avss.t116 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X264 multiplexer_0.trans_gate_m_32.in.t3 multiplexer_0.vtrip_1.t8 multiplexer_0.trans_gate_m_21.in.t3 avss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X265 avss.t143 avss.t144 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X266 a_n12118_9003# a_n8898_9381# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X267 avss.t96 avss.t97 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X268 a_n12654_n1203# a_n8898_n1203# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X269 multiplexer_0.trans_gate_m_29.in.t3 multiplexer_0.vtrip_0.t12 multiplexer_0.in_0011.t1 avss.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X270 dvdd.t32 dvdd.t29 dvdd.t31 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X271 multiplexer_0.in_1110.t2 multiplexer_0.in_1111.t2 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X272 dvdd.t28 dvdd.t25 dvdd.t27 dvdd.t26 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X273 a_n15874_5601# a_n12654_5223# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X274 multiplexer_0.vtrip_2_b.t0 multiplexer_0.vtrip_2.t5 avdd.t10 avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X275 a_n15874_2577# a_n12654_2955# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X276 multiplexer_0.trans_gate_m_21.in.t2 multiplexer_0.vtrip_0_b.t12 multiplexer_0.in_1011.t3 avdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X277 a_n8898_n1959# a_n5142_n1959.t1 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X278 dvdd.t24 dvdd.t22 dvdd.t23 dvdd.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X279 avss.t225 avss.t226 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X280 a_n12118_12783# a_n8898_12405# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X281 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.vtrip_0_b.t13 multiplexer_0.in_1100.t2 avss.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X282 dvss.t5 vtrip[3].t3 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X283 a_n8362_7869# multiplexer_0.in_0001.t2 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X284 a_n15874_13161# a_n12654_12783# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X285 comp_hyst_0.net3.t1 comp_hyst_0.net3.t0 dvdd.t101 dvdd.t26 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X286 ovout.t0 comp_hyst_0.net3.t0 dvdd.t100 dvdd.t99 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
X287 a_n12654_n447# a_n8898_n447# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X288 avss.t165 avss.t166 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X289 dvdd.t21 dvdd.t18 dvdd.t20 dvdd.t19 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X290 a_n8362_11649# a_n5142_12027# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X291 avss.t250 multiplexer_0.vtrip_3.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X292 avss.t77 avss.t78 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X293 a_n12118_9003# a_n8898_8625# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X294 a_n12118_5979# a_n8898_6357# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X295 dvdd.t17 dvdd.t14 dvdd.t16 dvdd.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X296 avss.t137 avss.t138 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X297 multiplexer_0.trans_gate_m_25.in.t1 multiplexer_0.vtrip_0.t13 multiplexer_0.in_0111.t1 avss.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X298 dvdd.t13 dvdd.t11 dvdd.t12 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X299 a_n15874_n1203# a_n12654_n825# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X300 avss.t212 avss.t213 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X301 a_n12118_12027# a_n8898_12405# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X302 avss.t32 avss.t33 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X303 comp_hyst_0.net4 comp_hyst_0.net3.t0 dvdd.t98 dvdd.t15 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X304 avss.t163 avss.t164 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X305 multiplexer_0.in_0101.t0 multiplexer_0.in_0110.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X306 avss.t75 avss.t76 avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X307 a_n15874_10137# a_n12654_9759# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X308 level_shifter_0.out multiplexer_0.vtrip_0_b.t14 avdd.t25 avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X309 multiplexer_0.in_1100.t0 multiplexer_0.in_1011.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X310 a_n15874_6357# a_n12654_6735# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X311 multiplexer_0.trans_gate_m_27.in.t3 multiplexer_0.vtrip_0_b.t15 multiplexer_0.in_0101.t3 avdd.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X312 avss.t206 avss.t207 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X313 avss.t132 vtrip[2].t2 multiplexer_0.vtrip_2_b.t1 avss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X314 a_n12118_3711# a_n8898_3333# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X315 dvss.t55 dvss.t53 dvss.t54 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X316 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.vtrip_0_b.t16 multiplexer_0.in_0000.t2 avss.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X317 avss.t204 avss.t205 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X318 a_n15874_13917# a_n12654_14295# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X319 vin.t0 multiplexer_0.vtrip_3.t5 multiplexer_0.trans_gate_m_33.in.t4 avdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X320 avss.t200 avss.t201 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X321 a_n15874_13917# a_n12654_13539# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X322 avss.t198 avss.t199 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X323 avss.t196 avss.t197 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X324 multiplexer_0.trans_gate_m_37.out.t3 multiplexer_0.vtrip_2.t6 multiplexer_0.trans_gate_m_37.in.t1 avss.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X325 dvss.t6 vin.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X326 a_n8362_10893# a_n5142_10515# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X327 a_n8898_687# a_n5142_687# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X328 avss.t194 avss.t195 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X329 avss.t257 avss.t258 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X330 a_n15874_4089# a_n12654_3711# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X331 multiplexer_0.trans_gate_m_19.in.t0 multiplexer_0.vtrip_0.t14 multiplexer_0.in_1110.t0 avdd.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X332 avss.t13 multiplexer_0.vtrip_2_b.t6 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X333 comp_hyst_0.net4 comp_hyst_0.net4 dvdd.t114 dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X334 a_n8898_n825# a_n5142_n825# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X335 comp_hyst_0.net3.t3 ena.t7 dvdd.t95 dvdd.t94 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X336 a_n12118_13539# a_n8898_13161# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X337 a_n12654_1065# a_n8898_1065# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X338 avss.t192 avss.t193 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X339 multiplexer_0.trans_gate_m_31.out.t2 multiplexer_0.vtrip_1_b.t10 multiplexer_0.trans_gate_m_31.in.t5 avss.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X340 multiplexer_0.trans_gate_m_37.in.t1 multiplexer_0.vtrip_1_b.t11 multiplexer_0.trans_gate_m_18.in.t5 avss.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X341 multiplexer_0.in_0100.t0 multiplexer_0.in_0011.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X342 avss.t50 avss.t51 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X343 comp_hyst_0.net3.t0 comp_hyst_0.net4 dvdd.t113 dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X344 avss.t135 avss.t136 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X345 a_n15874_7869# a_n12654_7491# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X346 avss.t93 avss.t94 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X347 dvss.t52 dvss.t50 dvss.t51 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X348 a_n15874_n1959# a_n12654_n1581# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X349 a_n8362_10137# a_n5142_10515# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X350 dvss.t17 vtrip[0].t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X351 multiplexer_0.trans_gate_m_33.in.t1 multiplexer_0.vtrip_2_b.t7 multiplexer_0.trans_gate_m_28.in.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X352 avss.t131 multiplexer_0.vtrip_0_b.t17 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X353 a_n8898_309# a_n5142_n69# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X354 avss.t234 avss.t235 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X355 a_n12118_4467# a_n8898_4845# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X356 avss.t11 avss.t12 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X357 dvss.t3 comp_hyst_0.net5 comp_hyst_0.net5.t0 dvss.t2 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X358 a_n15874_1065# a_n12654_1443# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X359 a_n12118_11271# a_n8898_10893# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X360 dvss.t49 dvss.t47 dvss.t48 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X361 avss.t232 avss.t233 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X362 a_n8898_14673# a_n5142_14295# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X363 dvss.t73 comp_hyst_0.net2 ovout.t2 dvss.t72 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
X364 multiplexer_0.in_1000.t3 multiplexer_0.in_1001.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X365 dvss.t19 vtrip[0].t3 level_shifter_0.in_b.t1 dvss.t18 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X366 dvss.t71 comp_hyst_0.ena_b.t1 ovout.t1 dvss.t70 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X367 avss.t148 avss.t149 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X368 multiplexer_0.trans_gate_m_28.in.t3 multiplexer_0.vtrip_1_b.t12 multiplexer_0.trans_gate_m_25.in.t5 avdd.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X369 avss.t73 avss.t74 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X370 a_n15874_n1203# a_n12654_n1203# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X371 multiplexer_0.trans_gate_m_21.in.t5 multiplexer_0.vtrip_0_b.t18 multiplexer_0.in_1010.t3 avss.t219 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X372 a_n12118_2199# a_n8898_1821# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X373 avss.t113 avss.t114 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X374 avss.t70 avss.t71 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X375 dvss.t46 dvss.t44 dvss.t45 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X376 a_n8362_7869# multiplexer_0.in_0010.t0 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X377 a_n15874_12405# a_n12654_12783# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X378 avss.t52 avss.t53 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X379 avss.t236 avss.t237 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X380 avss.t185 multiplexer_0.vtrip_1.t9 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X381 dvdd.t10 dvdd.t8 dvdd.t9 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X382 multiplexer_0.trans_gate_m_25.in.t0 multiplexer_0.vtrip_0.t15 multiplexer_0.in_0110.t2 avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X383 avss.t251 avss.t252 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X384 avss.t21 avss.t22 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X385 dvss.t43 dvss.t41 dvss.t42 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X386 multiplexer_0.trans_gate_m_23.in.t0 multiplexer_0.vtrip_0.t16 multiplexer_0.in_1000.t1 avdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X387 a_n8362_11649# a_n5142_11271# avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X388 a_n12118_8247# a_n8898_8625# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X389 a_n8898_1443# multiplexer_0.in_1111.t3 avss.t1 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X390 dvss.t40 dvss.t38 dvss.t39 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X391 a_n15874_4845# a_n12654_5223# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X392 multiplexer_0.vtrip_1_b.t1 level_shifter_1.out avdd.t29 avdd.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X393 dvss.t37 dvss.t35 dvss.t36 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X394 a_n12118_5979# a_n8898_5601# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X395 a_n15874_2577# a_n12654_2199# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X396 a_n12654_15051# a_n8898_15051# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X397 dvdd.t7 dvdd.t4 dvdd.t6 dvdd.t5 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X398 multiplexer_0.trans_gate_m_31.in.t0 multiplexer_0.vtrip_0.t17 multiplexer_0.in_0001.t1 avss.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X399 vin.t2 multiplexer_0.vtrip_3_b.t5 multiplexer_0.trans_gate_m_37.out.t5 avdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X400 dvss.t34 dvss.t32 dvss.t33 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X401 dvss.t31 dvss.t28 dvss.t30 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X402 ibias.t0 comp_hyst_0.ena_b comp_hyst_0.net5.t1 dvdd.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=5
X403 a_n15874_9381# a_n12654_9003# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X404 a_n15874_12405# a_n12654_12027# avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X405 a_n12654_n1959# a_n8898_n1959# avss.t2 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X406 dvss.t27 dvss.t24 dvss.t26 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X407 avss.t208 avss.t209 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X408 multiplexer_0.trans_gate_m_19.in.t3 multiplexer_0.vtrip_0_b.t19 multiplexer_0.in_1111.t1 avdd.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X409 multiplexer_0.trans_gate_m_27.in.t2 multiplexer_0.vtrip_0_b.t20 multiplexer_0.in_0100.t2 avss.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X410 avss.t238 avss.t239 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X411 avss.t4 avss.t5 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X412 avss.t48 avss.t49 avss.t3 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X413 dvdd.t3 dvdd.t0 dvdd.t2 dvdd.t1 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X414 avss.t174 avss.t175 avss.t8 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X415 dvss.t23 vtrip[2].t3 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
R0 dvss.n449 dvss.n444 254820
R1 dvss.n95 dvss.n94 34996.5
R2 dvss.n94 dvss.n9 31135.3
R3 dvss.n448 dvss.n447 30031.7
R4 dvss.n449 dvss.n448 23444.7
R5 dvss.n533 dvss.n21 17898.5
R6 dvss.n447 dvss.n444 14868.9
R7 dvss.n510 dvss.n54 13807.4
R8 dvss.n510 dvss.n50 13807.4
R9 dvss.n277 dvss.n49 13807.4
R10 dvss.n513 dvss.n49 13807.4
R11 dvss.n566 dvss.n9 13404.2
R12 dvss.n511 dvss.n51 12416.8
R13 dvss.n512 dvss.n511 12416.8
R14 dvss.n464 dvss.n10 11008.6
R15 dvss.n565 dvss.n10 11008.6
R16 dvss.n566 dvss.n565 11008.6
R17 dvss.n528 dvss.n40 6854.44
R18 dvss.n528 dvss.n41 6854.44
R19 dvss.n73 dvss.n41 6854.44
R20 dvss.n73 dvss.n40 6854.44
R21 dvss.n94 dvss.n93 6401.06
R22 dvss.n450 dvss.n443 4698.47
R23 dvss.t20 dvss.n113 4082.08
R24 dvss.n227 dvss.n114 4040.64
R25 dvss.n114 dvss.n105 4040.64
R26 dvss.n250 dvss.n96 4040.64
R27 dvss.n237 dvss.n96 4040.64
R28 dvss.n305 dvss.n69 3957.38
R29 dvss.n302 dvss.n69 3957.38
R30 dvss.n305 dvss.n70 3957.38
R31 dvss.n302 dvss.n70 3957.38
R32 dvss.n460 dvss.n457 3957.38
R33 dvss.n469 dvss.n457 3957.38
R34 dvss.n460 dvss.n459 3957.38
R35 dvss.n484 dvss.n481 3957.38
R36 dvss.n492 dvss.n481 3957.38
R37 dvss.n484 dvss.n483 3957.38
R38 dvss.n552 dvss.n16 3957.38
R39 dvss.n556 dvss.n16 3957.38
R40 dvss.n552 dvss.n18 3957.38
R41 dvss.n299 dvss.n283 3957.38
R42 dvss.n299 dvss.n297 3957.38
R43 dvss.n520 dvss.n516 3957.38
R44 dvss.n521 dvss.n520 3957.38
R45 dvss.n531 dvss.n37 3957.38
R46 dvss.n37 dvss.n35 3957.38
R47 dvss.n36 dvss.n35 3957.38
R48 dvss.n548 dvss.n5 3957.38
R49 dvss.n548 dvss.n546 3957.38
R50 dvss.n571 dvss.n5 3957.38
R51 dvss.n251 dvss.n95 3484.39
R52 dvss.n309 dvss.n308 3186.08
R53 dvss.n127 dvss.n116 3171.26
R54 dvss.n116 dvss.n115 3171.26
R55 dvss.n240 dvss.n112 3171.26
R56 dvss.n240 dvss.n107 3171.26
R57 dvss.n125 dvss.n117 3171.26
R58 dvss.n117 dvss.n106 3171.26
R59 dvss.n124 dvss.n118 3171.26
R60 dvss.n118 dvss.n101 3171.26
R61 dvss.n239 dvss.n238 3171.26
R62 dvss.n239 dvss.n97 3171.26
R63 dvss.n537 dvss.n27 3052.71
R64 dvss.n537 dvss.n536 3052.71
R65 dvss.n536 dvss.n535 3052.71
R66 dvss.n535 dvss.n27 3052.71
R67 dvss.n550 dvss.n21 2973.47
R68 dvss.n446 dvss.n443 2848.04
R69 dvss.n291 dvss.n283 2566.79
R70 dvss.n291 dvss.n290 2566.79
R71 dvss.n290 dvss.n42 2566.79
R72 dvss.n516 dvss.n42 2566.79
R73 dvss.n297 dvss.n284 2566.79
R74 dvss.n289 dvss.n284 2566.79
R75 dvss.n289 dvss.n43 2566.79
R76 dvss.n521 dvss.n43 2566.79
R77 dvss.n21 dvss.n9 2126.29
R78 dvss.n459 dvss.n455 1836.74
R79 dvss.n483 dvss.n479 1836.74
R80 dvss.n18 dvss.n15 1836.74
R81 dvss.n546 dvss.n3 1836.74
R82 dvss.n84 dvss.n58 1735.47
R83 dvss.n312 dvss.n58 1735.47
R84 dvss.n253 dvss.n92 1735.47
R85 dvss.n187 dvss.n181 1735.47
R86 dvss.n187 dvss.n157 1735.47
R87 dvss.n171 dvss.n170 1735.47
R88 dvss.n465 dvss.n458 1720.85
R89 dvss.n488 dvss.n482 1720.85
R90 dvss.n564 dvss.n11 1720.85
R91 dvss.n567 dvss.n6 1720.85
R92 dvss.t0 dvss.n19 1584.72
R93 dvss.n465 dvss.n456 1552.82
R94 dvss.n472 dvss.n456 1552.82
R95 dvss.n488 dvss.n480 1552.82
R96 dvss.n495 dvss.n480 1552.82
R97 dvss.n564 dvss.n12 1552.82
R98 dvss.n559 dvss.n12 1552.82
R99 dvss.n540 dvss.n22 1552.82
R100 dvss.n544 dvss.n22 1552.82
R101 dvss.n540 dvss.n23 1552.82
R102 dvss.n544 dvss.n23 1552.82
R103 dvss.n149 dvss.n132 1552.82
R104 dvss.n133 dvss.n132 1552.82
R105 dvss.n149 dvss.n148 1552.82
R106 dvss.n148 dvss.n133 1552.82
R107 dvss.n220 dvss.n219 1552.82
R108 dvss.n221 dvss.n220 1552.82
R109 dvss.n222 dvss.n219 1552.82
R110 dvss.n222 dvss.n221 1552.82
R111 dvss.n574 dvss.n4 1552.82
R112 dvss.n567 dvss.n4 1552.82
R113 dvss.n469 dvss.n458 1390.59
R114 dvss.n492 dvss.n482 1390.59
R115 dvss.n556 dvss.n11 1390.59
R116 dvss.n525 dvss.n42 1390.59
R117 dvss.n525 dvss.n43 1390.59
R118 dvss.n292 dvss.n291 1390.59
R119 dvss.n292 dvss.n284 1390.59
R120 dvss.n54 dvss.n51 1390.59
R121 dvss.n277 dvss.n51 1390.59
R122 dvss.n513 dvss.n512 1390.59
R123 dvss.n512 dvss.n50 1390.59
R124 dvss.n571 dvss.n6 1390.59
R125 dvss.t21 dvss.n20 1254.31
R126 dvss.n551 dvss.t8 1254.31
R127 dvss.n549 dvss.t18 1254.31
R128 dvss.n471 dvss.t0 1133.98
R129 dvss.n169 dvss.t25 1114.84
R130 dvss.n252 dvss.t29 1114.84
R131 dvss.n271 dvss.n60 968.173
R132 dvss.n60 dvss.n57 968.173
R133 dvss.n259 dvss.n79 968.173
R134 dvss.n270 dvss.n79 968.173
R135 dvss.n270 dvss.n269 968.173
R136 dvss.n269 dvss.n80 968.173
R137 dvss.n64 dvss.n59 968.173
R138 dvss.n260 dvss.n59 968.173
R139 dvss.n260 dvss.n62 968.173
R140 dvss.n271 dvss.n62 968.173
R141 dvss.n267 dvss.n85 968.173
R142 dvss.n267 dvss.n87 968.173
R143 dvss.n87 dvss.n82 968.173
R144 dvss.n259 dvss.n82 968.173
R145 dvss.n310 dvss.n63 968.173
R146 dvss.n310 dvss.n64 968.173
R147 dvss.n107 dvss.n104 968.173
R148 dvss.n115 dvss.n104 968.173
R149 dvss.n229 dvss.n125 968.173
R150 dvss.n229 dvss.n112 968.173
R151 dvss.n126 dvss.n112 968.173
R152 dvss.n127 dvss.n126 968.173
R153 dvss.n103 dvss.n101 968.173
R154 dvss.n106 dvss.n103 968.173
R155 dvss.n244 dvss.n106 968.173
R156 dvss.n244 dvss.n107 968.173
R157 dvss.n238 dvss.n120 968.173
R158 dvss.n124 dvss.n120 968.173
R159 dvss.n231 dvss.n124 968.173
R160 dvss.n231 dvss.n125 968.173
R161 dvss.n246 dvss.n97 968.173
R162 dvss.n246 dvss.n101 968.173
R163 dvss.n203 dvss.n156 968.173
R164 dvss.n192 dvss.n156 968.173
R165 dvss.n208 dvss.n178 968.173
R166 dvss.n208 dvss.n182 968.173
R167 dvss.n182 dvss.n180 968.173
R168 dvss.n191 dvss.n180 968.173
R169 dvss.n160 dvss.n155 968.173
R170 dvss.n197 dvss.n155 968.173
R171 dvss.n197 dvss.n158 968.173
R172 dvss.n203 dvss.n158 968.173
R173 dvss.n177 dvss.n164 968.173
R174 dvss.n211 dvss.n177 968.173
R175 dvss.n211 dvss.n210 968.173
R176 dvss.n210 dvss.n178 968.173
R177 dvss.n216 dvss.n159 968.173
R178 dvss.n216 dvss.n160 968.173
R179 dvss.n494 dvss.t21 897.556
R180 dvss.n558 dvss.t8 897.556
R181 dvss.n573 dvss.t18 897.556
R182 dvss.n84 dvss.n80 869.38
R183 dvss.n312 dvss.n57 869.38
R184 dvss.n90 dvss.n63 869.38
R185 dvss.n253 dvss.n85 869.38
R186 dvss.n227 dvss.n127 869.38
R187 dvss.n115 dvss.n105 869.38
R188 dvss.n250 dvss.n97 869.38
R189 dvss.n238 dvss.n237 869.38
R190 dvss.n191 dvss.n181 869.38
R191 dvss.n192 dvss.n157 869.38
R192 dvss.n170 dvss.n159 869.38
R193 dvss.n173 dvss.n164 869.38
R194 dvss.n139 dvss.n80 866.087
R195 dvss.n139 dvss.n57 866.087
R196 dvss.n272 dvss.n270 866.087
R197 dvss.n272 dvss.n271 866.087
R198 dvss.n261 dvss.n259 866.087
R199 dvss.n261 dvss.n260 866.087
R200 dvss.n87 dvss.n86 866.087
R201 dvss.n86 dvss.n64 866.087
R202 dvss.n255 dvss.n85 866.087
R203 dvss.n255 dvss.n63 866.087
R204 dvss.n193 dvss.n191 866.087
R205 dvss.n193 dvss.n192 866.087
R206 dvss.n204 dvss.n182 866.087
R207 dvss.n204 dvss.n203 866.087
R208 dvss.n198 dvss.n178 866.087
R209 dvss.n198 dvss.n197 866.087
R210 dvss.n212 dvss.n211 866.087
R211 dvss.n212 dvss.n160 866.087
R212 dvss.n165 dvss.n164 866.087
R213 dvss.n165 dvss.n159 866.087
R214 dvss.n275 dvss.n52 800.378
R215 dvss.n52 dvss.n48 800.378
R216 dvss.n458 dvss.n455 730.059
R217 dvss.n482 dvss.n479 730.059
R218 dvss.n15 dvss.n11 730.059
R219 dvss.n6 dvss.n3 730.059
R220 dvss.n91 dvss.n90 686.495
R221 dvss.n173 dvss.n172 686.495
R222 dvss.n472 dvss.n455 654.736
R223 dvss.n495 dvss.n479 654.736
R224 dvss.n559 dvss.n15 654.736
R225 dvss.n574 dvss.n3 654.736
R226 dvss.n543 dvss.n542 627.953
R227 dvss.n464 dvss.t5 543.74
R228 dvss.n169 dvss.n113 474.76
R229 dvss.n252 dvss.n251 474.76
R230 dvss.n249 dvss.n98 466.447
R231 dvss.n236 dvss.n98 466.447
R232 dvss.n471 dvss.n470 450.733
R233 dvss.n74 dvss.n72 445.365
R234 dvss.t23 dvss.n10 430.373
R235 dvss.n565 dvss.t7 430.373
R236 dvss.n566 dvss.t17 430.373
R237 dvss.n542 dvss.n541 429.183
R238 dvss.t20 dvss.n119 396.166
R239 dvss.n534 dvss.t16 374.048
R240 dvss.n538 dvss.t16 374.048
R241 dvss.n235 dvss.n99 362.541
R242 dvss.n248 dvss.n99 362.541
R243 dvss.n233 dvss.n121 362.541
R244 dvss.n121 dvss.n100 362.541
R245 dvss.n123 dvss.n122 362.541
R246 dvss.n122 dvss.n109 362.541
R247 dvss.n241 dvss.n111 362.541
R248 dvss.n242 dvss.n241 362.541
R249 dvss.n134 dvss.n129 362.541
R250 dvss.n135 dvss.n134 362.541
R251 dvss.n494 dvss.n493 356.757
R252 dvss.n558 dvss.n557 356.757
R253 dvss.n573 dvss.n572 356.757
R254 dvss.n30 dvss.n29 353.507
R255 dvss.n72 dvss.n38 348.613
R256 dvss.n102 dvss.n95 331.055
R257 dvss.n451 dvss.n442 305.281
R258 dvss.n465 dvss.n464 303.233
R259 dvss.n488 dvss.n10 300.995
R260 dvss.n565 dvss.n564 300.995
R261 dvss.n567 dvss.n566 300.995
R262 dvss.n542 dvss.n23 293.281
R263 dvss.n466 dvss.n465 292.5
R264 dvss.n463 dvss.n456 292.5
R265 dvss.t5 dvss.n456 292.5
R266 dvss.n473 dvss.n472 292.5
R267 dvss.n472 dvss.n471 292.5
R268 dvss.n489 dvss.n488 292.5
R269 dvss.n487 dvss.n480 292.5
R270 dvss.t23 dvss.n480 292.5
R271 dvss.n496 dvss.n495 292.5
R272 dvss.n495 dvss.n494 292.5
R273 dvss.n564 dvss.n563 292.5
R274 dvss.n562 dvss.n12 292.5
R275 dvss.n12 dvss.t7 292.5
R276 dvss.n560 dvss.n559 292.5
R277 dvss.n559 dvss.n558 292.5
R278 dvss.n221 dvss.n152 292.5
R279 dvss.n221 dvss.n119 292.5
R280 dvss.n223 dvss.n222 292.5
R281 dvss.n222 dvss.t6 292.5
R282 dvss.n219 dvss.n154 292.5
R283 dvss.n219 dvss.n218 292.5
R284 dvss.n220 dvss.n130 292.5
R285 dvss.n220 dvss.t6 292.5
R286 dvss.n145 dvss.n133 292.5
R287 dvss.n133 dvss.n83 292.5
R288 dvss.n148 dvss.n147 292.5
R289 dvss.n148 dvss.t10 292.5
R290 dvss.n150 dvss.n149 292.5
R291 dvss.n149 dvss.n102 292.5
R292 dvss.n138 dvss.n132 292.5
R293 dvss.n132 dvss.t10 292.5
R294 dvss.n544 dvss.n543 292.5
R295 dvss.n545 dvss.n544 292.5
R296 dvss.n23 dvss.t11 292.5
R297 dvss.n541 dvss.n540 292.5
R298 dvss.n540 dvss.n539 292.5
R299 dvss.n24 dvss.n22 292.5
R300 dvss.n22 dvss.t11 292.5
R301 dvss.n8 dvss.n4 292.5
R302 dvss.t17 dvss.n4 292.5
R303 dvss.n568 dvss.n567 292.5
R304 dvss.n575 dvss.n574 292.5
R305 dvss.n574 dvss.n573 292.5
R306 dvss.n515 dvss.n47 292.142
R307 dvss.n515 dvss.n514 292.142
R308 dvss.n462 dvss.n461 257.13
R309 dvss.n486 dvss.n485 257.13
R310 dvss.n554 dvss.n553 257.13
R311 dvss.n47 dvss.n46 257.13
R312 dvss.n547 dvss.n7 257.13
R313 dvss.n29 dvss.n28 246.004
R314 dvss.n570 dvss.n7 215.569
R315 dvss.n303 dvss.n71 215.506
R316 dvss.n533 dvss.t14 215.23
R317 dvss.n298 dvss.t70 203.126
R318 dvss.t68 dvss.n53 203.126
R319 dvss.n526 dvss.t12 203.126
R320 dvss.n89 dvss.n88 202.918
R321 dvss.n254 dvss.n88 202.918
R322 dvss.n168 dvss.n167 202.918
R323 dvss.n174 dvss.n167 202.918
R324 dvss.n533 dvss.n31 192.123
R325 dvss.n550 dvss.n19 189.595
R326 dvss.n445 dvss.n442 185.155
R327 dvss.n468 dvss.n462 175.536
R328 dvss.n491 dvss.n486 175.536
R329 dvss.n555 dvss.n554 175.536
R330 dvss.t70 dvss.t74 173.322
R331 dvss.n46 dvss.n38 169.59
R332 dvss.t14 dvss.t12 160.484
R333 dvss.n33 dvss.n31 160.484
R334 dvss.n311 dvss.n61 150.856
R335 dvss.n550 dvss.n20 150.065
R336 dvss.n551 dvss.n550 150.065
R337 dvss.n550 dvss.n549 150.065
R338 dvss.n316 dvss.n30 148.329
R339 dvss.n527 dvss.n34 146.728
R340 dvss.n550 dvss.n545 129.994
R341 dvss.n315 dvss.n50 126.078
R342 dvss.n414 dvss.t38 125.236
R343 dvss.t38 dvss.n413 125.236
R344 dvss.n394 dvss.t62 125.236
R345 dvss.t62 dvss.n393 125.236
R346 dvss.n390 dvss.t65 125.236
R347 dvss.t65 dvss.n389 125.236
R348 dvss.n386 dvss.t35 125.236
R349 dvss.t35 dvss.n385 125.236
R350 dvss.n382 dvss.t24 125.236
R351 dvss.t24 dvss.n381 125.236
R352 dvss.t41 dvss.n417 125.236
R353 dvss.n418 dvss.t41 125.236
R354 dvss.n323 dvss.t47 125.236
R355 dvss.t47 dvss.n322 125.236
R356 dvss.n321 dvss.t44 125.236
R357 dvss.t44 dvss.n320 125.236
R358 dvss.n445 dvss.n444 122.587
R359 dvss.n209 dvss.t25 120.593
R360 dvss.n311 dvss.t29 120.593
R361 dvss.n316 dvss.n25 120.013
R362 dvss.n373 dvss.t53 118.005
R363 dvss.t53 dvss.n372 118.005
R364 dvss.n360 dvss.t50 118.005
R365 dvss.t50 dvss.n355 118.005
R366 dvss.n410 dvss.t28 118.005
R367 dvss.t28 dvss.n409 118.005
R368 dvss.n400 dvss.t59 118.005
R369 dvss.t59 dvss.n399 118.005
R370 dvss.n469 dvss.n468 117.001
R371 dvss.n470 dvss.n469 117.001
R372 dvss.n461 dvss.n460 117.001
R373 dvss.n460 dvss.n19 117.001
R374 dvss.n492 dvss.n491 117.001
R375 dvss.n493 dvss.n492 117.001
R376 dvss.n485 dvss.n484 117.001
R377 dvss.n484 dvss.n20 117.001
R378 dvss.n556 dvss.n555 117.001
R379 dvss.n557 dvss.n556 117.001
R380 dvss.n553 dvss.n552 117.001
R381 dvss.n552 dvss.n551 117.001
R382 dvss.n171 dvss.n167 117.001
R383 dvss.n166 dvss.n165 117.001
R384 dvss.n165 dvss.t25 117.001
R385 dvss.n92 dvss.n88 117.001
R386 dvss.n256 dvss.n255 117.001
R387 dvss.n255 dvss.t29 117.001
R388 dvss.n47 dvss.n35 117.001
R389 dvss.t14 dvss.n35 117.001
R390 dvss.n531 dvss.n530 117.001
R391 dvss.n213 dvss.n212 117.001
R392 dvss.n212 dvss.t25 117.001
R393 dvss.n199 dvss.n198 117.001
R394 dvss.n198 dvss.t25 117.001
R395 dvss.n205 dvss.n204 117.001
R396 dvss.n204 dvss.t25 117.001
R397 dvss.n194 dvss.n193 117.001
R398 dvss.n193 dvss.t25 117.001
R399 dvss.n188 dvss.n187 117.001
R400 dvss.n187 dvss.t25 117.001
R401 dvss.n514 dvss.n513 117.001
R402 dvss.n513 dvss.n31 117.001
R403 dvss.n50 dvss.n31 117.001
R404 dvss.n55 dvss.n54 117.001
R405 dvss.n61 dvss.n54 117.001
R406 dvss.n278 dvss.n277 117.001
R407 dvss.n277 dvss.n61 117.001
R408 dvss.n293 dvss.n292 117.001
R409 dvss.n292 dvss.n53 117.001
R410 dvss.n525 dvss.n524 117.001
R411 dvss.n526 dvss.n525 117.001
R412 dvss.n520 dvss.n519 117.001
R413 dvss.n520 dvss.n33 117.001
R414 dvss.n300 dvss.n299 117.001
R415 dvss.n299 dvss.n298 117.001
R416 dvss.n281 dvss.n70 117.001
R417 dvss.t72 dvss.n70 117.001
R418 dvss.n69 dvss.n66 117.001
R419 dvss.t72 dvss.n69 117.001
R420 dvss.n529 dvss.n528 117.001
R421 dvss.n528 dvss.n527 117.001
R422 dvss.n74 dvss.n73 117.001
R423 dvss.n73 dvss.n71 117.001
R424 dvss.n86 dvss.n67 117.001
R425 dvss.n86 dvss.t29 117.001
R426 dvss.n262 dvss.n261 117.001
R427 dvss.n261 dvss.t29 117.001
R428 dvss.n273 dvss.n272 117.001
R429 dvss.n272 dvss.t29 117.001
R430 dvss.n140 dvss.n139 117.001
R431 dvss.n139 dvss.t29 117.001
R432 dvss.n144 dvss.n58 117.001
R433 dvss.t29 dvss.n58 117.001
R434 dvss.n571 dvss.n570 117.001
R435 dvss.n572 dvss.n571 117.001
R436 dvss.n548 dvss.n547 117.001
R437 dvss.n549 dvss.n548 117.001
R438 dvss.n235 dvss.n234 115.201
R439 dvss.n234 dvss.n233 115.201
R440 dvss.n248 dvss.n247 115.201
R441 dvss.n247 dvss.n100 115.201
R442 dvss.n108 dvss.n100 115.201
R443 dvss.n109 dvss.n108 115.201
R444 dvss.n233 dvss.n232 115.201
R445 dvss.n232 dvss.n123 115.201
R446 dvss.n228 dvss.n123 115.201
R447 dvss.n228 dvss.n111 115.201
R448 dvss.n243 dvss.n109 115.201
R449 dvss.n243 dvss.n242 115.201
R450 dvss.n242 dvss.n110 115.201
R451 dvss.n135 dvss.n110 115.201
R452 dvss.n128 dvss.n111 115.201
R453 dvss.n129 dvss.n128 115.201
R454 dvss.n81 dvss.n78 115.201
R455 dvss.n141 dvss.n81 115.201
R456 dvss.n263 dvss.n258 115.201
R457 dvss.n258 dvss.n78 115.201
R458 dvss.n265 dvss.n264 115.201
R459 dvss.n264 dvss.n263 115.201
R460 dvss.n266 dvss.n257 115.201
R461 dvss.n266 dvss.n265 115.201
R462 dvss.n309 dvss.n65 115.201
R463 dvss.n202 dvss.n196 115.201
R464 dvss.n196 dvss.n195 115.201
R465 dvss.n207 dvss.n183 115.201
R466 dvss.n207 dvss.n206 115.201
R467 dvss.n206 dvss.n184 115.201
R468 dvss.n190 dvss.n184 115.201
R469 dvss.n214 dvss.n162 115.201
R470 dvss.n200 dvss.n162 115.201
R471 dvss.n201 dvss.n200 115.201
R472 dvss.n202 dvss.n201 115.201
R473 dvss.n176 dvss.n175 115.201
R474 dvss.n176 dvss.n163 115.201
R475 dvss.n179 dvss.n163 115.201
R476 dvss.n183 dvss.n179 115.201
R477 dvss.n215 dvss.n161 115.201
R478 dvss.n215 dvss.n214 115.201
R479 dvss.n189 dvss.n188 112.451
R480 dvss.n532 dvss.n531 112.177
R481 dvss.n304 dvss.t72 111.421
R482 dvss.t72 dvss.n303 111.421
R483 dvss.n75 dvss.n66 104.514
R484 dvss.n249 dvss.n248 103.906
R485 dvss.n236 dvss.n235 103.906
R486 dvss.n226 dvss.n129 103.906
R487 dvss.n226 dvss.n225 103.906
R488 dvss.n136 dvss.n135 103.906
R489 dvss.n137 dvss.n136 103.906
R490 dvss.n142 dvss.n141 103.906
R491 dvss.n143 dvss.n142 103.906
R492 dvss.n89 dvss.n65 103.906
R493 dvss.n257 dvss.n254 103.906
R494 dvss.n190 dvss.n189 103.906
R495 dvss.n195 dvss.n186 103.906
R496 dvss.n186 dvss.n185 103.906
R497 dvss.n168 dvss.n161 103.906
R498 dvss.n175 dvss.n174 103.906
R499 dvss.n470 dvss.t5 103.74
R500 dvss.n461 dvss.n453 100.233
R501 dvss.n485 dvss.n477 100.233
R502 dvss.n553 dvss.n17 100.233
R503 dvss.n547 dvss.n1 100.233
R504 dvss.n141 dvss.n140 99.0123
R505 dvss.n273 dvss.n78 99.0123
R506 dvss.n263 dvss.n262 99.0123
R507 dvss.n265 dvss.n67 99.0123
R508 dvss.n257 dvss.n256 99.0123
R509 dvss.n256 dvss.n65 99.0123
R510 dvss.n194 dvss.n190 99.0123
R511 dvss.n195 dvss.n194 99.0123
R512 dvss.n206 dvss.n205 99.0123
R513 dvss.n205 dvss.n202 99.0123
R514 dvss.n199 dvss.n183 99.0123
R515 dvss.n200 dvss.n199 99.0123
R516 dvss.n213 dvss.n163 99.0123
R517 dvss.n214 dvss.n213 99.0123
R518 dvss.n175 dvss.n166 99.0123
R519 dvss.n166 dvss.n161 99.0123
R520 dvss.n174 dvss.n173 97.5005
R521 dvss.n170 dvss.n168 97.5005
R522 dvss.n170 dvss.n169 97.5005
R523 dvss.n237 dvss.n236 97.5005
R524 dvss.n237 dvss.n113 97.5005
R525 dvss.n250 dvss.n249 97.5005
R526 dvss.n251 dvss.n250 97.5005
R527 dvss.n254 dvss.n253 97.5005
R528 dvss.n253 dvss.n252 97.5005
R529 dvss.n90 dvss.n89 97.5005
R530 dvss.n189 dvss.n181 97.5005
R531 dvss.n209 dvss.n181 97.5005
R532 dvss.n186 dvss.n157 97.5005
R533 dvss.n217 dvss.n157 97.5005
R534 dvss.n227 dvss.n226 97.5005
R535 dvss.n230 dvss.n227 97.5005
R536 dvss.n136 dvss.n105 97.5005
R537 dvss.n245 dvss.n105 97.5005
R538 dvss.n142 dvss.n84 97.5005
R539 dvss.n268 dvss.n84 97.5005
R540 dvss.n313 dvss.n312 97.5005
R541 dvss.n312 dvss.n311 97.5005
R542 dvss.n535 dvss.n30 97.5005
R543 dvss.n535 dvss.n534 97.5005
R544 dvss.n537 dvss.n26 97.5005
R545 dvss.n538 dvss.n537 97.5005
R546 dvss.n514 dvss.n48 96.7534
R547 dvss.n524 dvss.n44 94.3698
R548 dvss.n140 dvss.n56 92.6123
R549 dvss.n276 dvss.n273 92.6123
R550 dvss.n262 dvss.n77 92.6123
R551 dvss.n307 dvss.n67 92.6123
R552 dvss.n304 dvss.n61 91.7054
R553 dvss.n524 dvss.n523 90.3534
R554 dvss.n293 dvss.n287 90.3534
R555 dvss.n294 dvss.n293 90.3534
R556 dvss.n308 dvss.n66 85.0829
R557 dvss.n423 dvss.t15 84.6474
R558 dvss.n422 dvss.t75 84.2828
R559 dvss.n476 dvss.t1 84.2462
R560 dvss.n499 dvss.t22 84.2462
R561 dvss.n501 dvss.t9 84.2462
R562 dvss.n0 dvss.t19 84.2462
R563 dvss.n318 dvss.t4 83.7172
R564 dvss.n429 dvss.t3 83.7172
R565 dvss.n420 dvss.t71 83.7172
R566 dvss.n425 dvss.t69 83.7172
R567 dvss.n421 dvss.t13 83.7172
R568 dvss.n177 dvss.n176 83.5719
R569 dvss.n209 dvss.n177 83.5719
R570 dvss.n216 dvss.n215 83.5719
R571 dvss.n217 dvss.n216 83.5719
R572 dvss.n210 dvss.n179 83.5719
R573 dvss.n210 dvss.n209 83.5719
R574 dvss.n162 dvss.n155 83.5719
R575 dvss.n217 dvss.n155 83.5719
R576 dvss.n208 dvss.n207 83.5719
R577 dvss.n209 dvss.n208 83.5719
R578 dvss.n201 dvss.n158 83.5719
R579 dvss.n217 dvss.n158 83.5719
R580 dvss.n184 dvss.n180 83.5719
R581 dvss.n209 dvss.n180 83.5719
R582 dvss.n196 dvss.n156 83.5719
R583 dvss.n217 dvss.n156 83.5719
R584 dvss.n234 dvss.n120 83.5719
R585 dvss.n230 dvss.n120 83.5719
R586 dvss.n247 dvss.n246 83.5719
R587 dvss.n246 dvss.n245 83.5719
R588 dvss.n232 dvss.n231 83.5719
R589 dvss.n231 dvss.n230 83.5719
R590 dvss.n108 dvss.n103 83.5719
R591 dvss.n245 dvss.n103 83.5719
R592 dvss.n229 dvss.n228 83.5719
R593 dvss.n230 dvss.n229 83.5719
R594 dvss.n244 dvss.n243 83.5719
R595 dvss.n245 dvss.n244 83.5719
R596 dvss.n128 dvss.n126 83.5719
R597 dvss.n230 dvss.n126 83.5719
R598 dvss.n110 dvss.n104 83.5719
R599 dvss.n245 dvss.n104 83.5719
R600 dvss.n267 dvss.n266 83.5719
R601 dvss.n268 dvss.n267 83.5719
R602 dvss.n310 dvss.n309 83.5719
R603 dvss.n311 dvss.n310 83.5719
R604 dvss.n264 dvss.n82 83.5719
R605 dvss.n268 dvss.n82 83.5719
R606 dvss.n68 dvss.n59 83.5719
R607 dvss.n311 dvss.n59 83.5719
R608 dvss.n258 dvss.n79 83.5719
R609 dvss.n268 dvss.n79 83.5719
R610 dvss.n279 dvss.n62 83.5719
R611 dvss.n311 dvss.n62 83.5719
R612 dvss.n269 dvss.n81 83.5719
R613 dvss.n269 dvss.n268 83.5719
R614 dvss.n274 dvss.n60 83.5719
R615 dvss.n311 dvss.n60 83.5719
R616 dvss.n438 dvss.t55 82.8472
R617 dvss.n359 dvss.t51 82.8472
R618 dvss.n354 dvss.t52 82.8472
R619 dvss.n364 dvss.t54 82.8472
R620 dvss.n407 dvss.t30 82.8472
R621 dvss.n397 dvss.t60 82.8472
R622 dvss.n332 dvss.t31 82.8472
R623 dvss.n334 dvss.t58 82.8472
R624 dvss.n336 dvss.t57 82.8472
R625 dvss.n338 dvss.t61 82.8472
R626 dvss.n363 dvss.t34 82.8472
R627 dvss.n356 dvss.t33 82.8472
R628 dvss.n493 dvss.t23 82.1112
R629 dvss.n557 dvss.t7 82.1112
R630 dvss.n572 dvss.t17 82.1112
R631 dvss.n433 dvss.t49 77.4826
R632 dvss.n436 dvss.t46 77.4826
R633 dvss.n369 dvss.t45 77.4826
R634 dvss.n366 dvss.t48 77.4826
R635 dvss.n326 dvss.t42 77.4826
R636 dvss.n324 dvss.t43 77.4826
R637 dvss.n330 dvss.t39 77.4826
R638 dvss.n328 dvss.t40 77.4826
R639 dvss.n339 dvss.t63 77.4826
R640 dvss.n344 dvss.t66 77.4826
R641 dvss.n348 dvss.t36 77.4826
R642 dvss.n352 dvss.t26 77.4826
R643 dvss.n350 dvss.t27 77.4826
R644 dvss.n346 dvss.t37 77.4826
R645 dvss.n342 dvss.t67 77.4826
R646 dvss.n341 dvss.t64 77.4826
R647 dvss.n569 dvss.n568 77.3462
R648 dvss.n569 dvss.n2 75.6711
R649 dvss.n83 dvss.t29 75.657
R650 dvss.n218 dvss.t25 75.1985
R651 dvss.n539 dvss.t11 73.3432
R652 dvss.n545 dvss.t11 73.3432
R653 dvss.n172 dvss.n171 66.2531
R654 dvss.n92 dvss.n91 66.2531
R655 dvss.t20 dvss.n95 58.3417
R656 dvss.n543 dvss.n24 57.3914
R657 dvss.n539 dvss.n538 56.418
R658 dvss.n298 dvss.n71 55.9405
R659 dvss.n534 dvss.n533 55.2896
R660 dvss.n459 dvss.n453 53.1823
R661 dvss.n459 dvss.t0 53.1823
R662 dvss.n462 dvss.n457 53.1823
R663 dvss.n457 dvss.t0 53.1823
R664 dvss.n483 dvss.n477 53.1823
R665 dvss.n483 dvss.t21 53.1823
R666 dvss.n486 dvss.n481 53.1823
R667 dvss.n481 dvss.t21 53.1823
R668 dvss.n18 dvss.n17 53.1823
R669 dvss.n18 dvss.t8 53.1823
R670 dvss.n554 dvss.n16 53.1823
R671 dvss.n16 dvss.t8 53.1823
R672 dvss.n46 dvss.n37 53.1823
R673 dvss.n93 dvss.n37 53.1823
R674 dvss.n522 dvss.n521 53.1823
R675 dvss.n521 dvss.t12 53.1823
R676 dvss.n289 dvss.n45 53.1823
R677 dvss.t68 dvss.n289 53.1823
R678 dvss.n297 dvss.n296 53.1823
R679 dvss.t70 dvss.n297 53.1823
R680 dvss.n285 dvss.n283 53.1823
R681 dvss.t70 dvss.n283 53.1823
R682 dvss.n290 dvss.n288 53.1823
R683 dvss.n290 dvss.t68 53.1823
R684 dvss.n517 dvss.n516 53.1823
R685 dvss.n516 dvss.t12 53.1823
R686 dvss.n302 dvss.n301 53.1823
R687 dvss.n303 dvss.n302 53.1823
R688 dvss.n306 dvss.n305 53.1823
R689 dvss.n305 dvss.n304 53.1823
R690 dvss.n518 dvss.n36 53.1823
R691 dvss.n7 dvss.n5 53.1823
R692 dvss.n5 dvss.t18 53.1823
R693 dvss.n546 dvss.n1 53.1823
R694 dvss.n546 dvss.t18 53.1823
R695 dvss.t68 dvss.n34 52.7308
R696 dvss.n147 dvss.n131 51.9534
R697 dvss.n147 dvss.n146 51.9534
R698 dvss.n223 dvss.n153 51.9534
R699 dvss.n224 dvss.n223 51.9534
R700 dvss.n532 dvss.n36 50.9901
R701 dvss.n466 dvss.n463 49.0248
R702 dvss.n489 dvss.n487 49.0248
R703 dvss.n563 dvss.n562 49.0248
R704 dvss.n568 dvss.n8 49.0248
R705 dvss.n172 dvss.t25 46.2824
R706 dvss.n91 dvss.t29 46.2824
R707 dvss.n75 dvss.n74 45.9798
R708 dvss.n245 dvss.n102 45.8529
R709 dvss.n218 dvss.n217 45.3944
R710 dvss.n230 dvss.n119 45.3944
R711 dvss.n268 dvss.n83 44.9359
R712 dvss.n93 dvss.n32 44.3777
R713 dvss.n467 dvss.n466 43.6573
R714 dvss.n490 dvss.n489 43.6573
R715 dvss.n563 dvss.n13 43.6573
R716 dvss.t14 dvss.n33 42.6433
R717 dvss.t74 dvss.n34 37.7211
R718 dvss.n315 dvss.n48 36.3262
R719 dvss.n467 dvss.n454 34.6358
R720 dvss.n490 dvss.n478 34.6358
R721 dvss.n561 dvss.n13 34.6358
R722 dvss.n29 dvss.n27 34.4123
R723 dvss.n27 dvss.t16 34.4123
R724 dvss.n536 dvss.n25 34.4123
R725 dvss.n536 dvss.t16 34.4123
R726 dvss.n522 dvss.n515 31.827
R727 dvss.n428 dvss.t73 30.767
R728 dvss.n509 dvss.n314 29.5006
R729 dvss.n152 dvss.n151 28.0695
R730 dvss.n151 dvss.n150 28.037
R731 dvss.n268 dvss.t10 26.1364
R732 dvss.n217 dvss.t6 25.6779
R733 dvss.n230 dvss.t6 25.6779
R734 dvss.n533 dvss.n32 25.5174
R735 dvss.n245 dvss.t10 25.2193
R736 dvss.n72 dvss.n40 23.4005
R737 dvss.n40 dvss.n32 23.4005
R738 dvss.n286 dvss.n41 23.4005
R739 dvss.t74 dvss.n41 23.4005
R740 dvss.n288 dvss.n287 23.0509
R741 dvss.n98 dvss.n96 22.5005
R742 dvss.t20 dvss.n96 22.5005
R743 dvss.n239 dvss.n99 22.5005
R744 dvss.t20 dvss.n239 22.5005
R745 dvss.n121 dvss.n118 22.5005
R746 dvss.t20 dvss.n118 22.5005
R747 dvss.n122 dvss.n117 22.5005
R748 dvss.t20 dvss.n117 22.5005
R749 dvss.n241 dvss.n240 22.5005
R750 dvss.n240 dvss.t20 22.5005
R751 dvss.n134 dvss.n116 22.5005
R752 dvss.t20 dvss.n116 22.5005
R753 dvss.n151 dvss.n114 22.5005
R754 dvss.t20 dvss.n114 22.5005
R755 dvss.n285 dvss.n76 22.1664
R756 dvss.n288 dvss.n44 21.7501
R757 dvss.n452 dvss.n451 21.6109
R758 dvss.t2 dvss.t74 20.1756
R759 dvss.n286 dvss.n285 19.6688
R760 dvss.n294 dvss.n45 18.5312
R761 dvss.n523 dvss.n45 18.5312
R762 dvss.n523 dvss.n522 18.5312
R763 dvss.n508 dvss.n317 18.0964
R764 dvss.n296 dvss.n282 17.8201
R765 dvss.n296 dvss.n295 17.6528
R766 dvss.n519 dvss.n518 17.4088
R767 dvss.n518 dvss.n517 15.6648
R768 dvss.n468 dvss.n467 15.1599
R769 dvss.n491 dvss.n490 15.1599
R770 dvss.n555 dvss.n13 15.1599
R771 dvss.n317 dvss.n315 14.2671
R772 dvss.n570 dvss.n569 14.1572
R773 dvss.n509 dvss.n508 13.7723
R774 dvss.n542 dvss.n25 13.1595
R775 dvss.n541 dvss.n26 12.8005
R776 dvss.t32 dvss.n376 11.7013
R777 dvss.n377 dvss.t32 11.7013
R778 dvss.t56 dvss.n404 11.7013
R779 dvss.n405 dvss.t56 11.7013
R780 dvss.n529 dvss.n39 11.2005
R781 dvss.n282 dvss.n281 10.4113
R782 dvss.n281 dvss.n280 10.1864
R783 dvss.t2 dvss.n53 9.62951
R784 dvss.n511 dvss.n52 9.59066
R785 dvss.n511 dvss.t2 9.59066
R786 dvss.n510 dvss.n509 9.59066
R787 dvss.t2 dvss.n510 9.59066
R788 dvss.n295 dvss.n49 9.59066
R789 dvss.t2 dvss.n49 9.59066
R790 dvss.n314 dvss.n55 8.46331
R791 dvss.n300 dvss.n282 8.03628
R792 dvss.n144 dvss.n56 7.99238
R793 dvss.n137 dvss.n131 7.92886
R794 dvss.n225 dvss.n224 7.83334
R795 dvss.n185 dvss.n153 7.83334
R796 dvss.n146 dvss.n143 7.73781
R797 dvss.n28 dvss.n24 7.52991
R798 dvss.n275 dvss.n274 7.47598
R799 dvss.n77 dvss.n68 7.34402
R800 dvss.n530 dvss.n38 7.08621
R801 dvss.n143 dvss.n138 6.74438
R802 dvss.t14 dvss.n34 6.65708
R803 dvss.n185 dvss.n130 6.61638
R804 dvss.n225 dvss.n130 6.61638
R805 dvss.n138 dvss.n137 6.48838
R806 dvss.n308 dvss.n307 6.25272
R807 dvss.n279 dvss.n278 6.24182
R808 dvss.n463 dvss.n454 5.62598
R809 dvss.n487 dvss.n478 5.62598
R810 dvss.n562 dvss.n561 5.62598
R811 dvss.n8 dvss.n2 5.62598
R812 dvss.n280 dvss.n279 5.45041
R813 dvss.n145 dvss.n144 5.36091
R814 dvss.n188 dvss.n154 5.32842
R815 dvss.n278 dvss.n276 5.14871
R816 dvss.n474 dvss.n473 4.81722
R817 dvss.n497 dvss.n496 4.81722
R818 dvss.n560 dvss.n14 4.81722
R819 dvss.n576 dvss.n575 4.81722
R820 dvss.n307 dvss.n306 4.13833
R821 dvss.n276 dvss.n275 3.91455
R822 dvss.n301 dvss.n76 3.78325
R823 dvss.n527 dvss.n526 3.6687
R824 dvss.n301 dvss.n300 3.64012
R825 dvss.n517 dvss.n39 3.4019
R826 dvss.n287 dvss.n286 3.38261
R827 dvss.n306 dvss.n68 3.20618
R828 dvss.n280 dvss.n77 2.68327
R829 dvss.n76 dvss.n75 2.51552
R830 dvss.n405 dvss.n335 2.25322
R831 dvss.n406 dvss.n405 2.25322
R832 dvss.n404 dvss.n402 2.25322
R833 dvss.n404 dvss.n403 2.25322
R834 dvss.n378 dvss.n377 2.25322
R835 dvss.n377 dvss.n357 2.25322
R836 dvss.n376 dvss.n362 2.25322
R837 dvss.n376 dvss.n375 2.25322
R838 dvss.n474 dvss.n453 2.25276
R839 dvss.n497 dvss.n477 2.25276
R840 dvss.n17 dvss.n14 2.25276
R841 dvss.n576 dvss.n1 2.25276
R842 dvss.n314 dvss.n313 2.11039
R843 dvss.n426 dvss.n421 1.86647
R844 dvss.n447 dvss.n446 1.70108
R845 dvss.n428 dvss.n427 1.60988
R846 dvss.n446 dvss.n445 1.59604
R847 dvss.n274 dvss.n55 1.58728
R848 dvss.t14 dvss.n532 1.50849
R849 dvss.n427 dvss.n426 1.38166
R850 dvss.n530 dvss.n529 1.30662
R851 dvss.n505 dvss.n504 1.23532
R852 dvss.n424 dvss.n422 1.2043
R853 dvss.n424 dvss.n423 1.2043
R854 dvss.n502 dvss.n0 1.08443
R855 dvss.n398 dvss.n335 1.03311
R856 dvss.n408 dvss.n406 1.03311
R857 dvss.n402 dvss.n401 1.03311
R858 dvss.n403 dvss.n333 1.03311
R859 dvss.n379 dvss.n378 1.03311
R860 dvss.n371 dvss.n357 1.03311
R861 dvss.n362 dvss.n361 1.03311
R862 dvss.n375 dvss.n374 1.03311
R863 dvss.n503 dvss.n502 0.979071
R864 dvss.n504 dvss.n503 0.978625
R865 dvss.n295 dvss.n294 0.878931
R866 dvss.n317 dvss.n316 0.780399
R867 dvss.n435 dvss.n434 0.7505
R868 dvss.n431 dvss.n430 0.714563
R869 dvss.n360 dvss.n359 0.709739
R870 dvss.n399 dvss.n397 0.709739
R871 dvss.n409 dvss.n332 0.709739
R872 dvss.n438 dvss.n437 0.688
R873 dvss.n429 dvss.n318 0.654856
R874 dvss.n44 dvss.n39 0.653561
R875 dvss.n358 dvss.n353 0.6255
R876 dvss.n380 dvss.n379 0.6255
R877 dvss.n351 dvss.n349 0.6255
R878 dvss.n384 dvss.n383 0.6255
R879 dvss.n347 dvss.n345 0.6255
R880 dvss.n388 dvss.n387 0.6255
R881 dvss.n343 dvss.n340 0.6255
R882 dvss.n392 dvss.n391 0.6255
R883 dvss.n396 dvss.n395 0.6255
R884 dvss.n401 dvss.n337 0.6255
R885 dvss.n333 dvss.n331 0.6255
R886 dvss.n412 dvss.n411 0.6255
R887 dvss.n329 dvss.n327 0.6255
R888 dvss.n416 dvss.n415 0.6255
R889 dvss.n365 dvss.n325 0.6255
R890 dvss.n368 dvss.n367 0.6255
R891 dvss.n371 dvss.n370 0.6255
R892 dvss.n439 dvss.n438 0.589954
R893 dvss.n431 dvss.n419 0.568435
R894 dvss.n507 dvss.n506 0.563319
R895 dvss.n146 dvss.n145 0.552784
R896 dvss.n224 dvss.n152 0.552784
R897 dvss.n150 dvss.n131 0.552784
R898 dvss.n154 dvss.n153 0.552784
R899 dvss.n430 dvss.n429 0.539326
R900 dvss.n440 dvss.n25 0.517167
R901 dvss.n433 dvss.n432 0.503217
R902 dvss.n434 dvss.n433 0.503217
R903 dvss.n436 dvss.n435 0.503217
R904 dvss.n437 dvss.n436 0.503217
R905 dvss.n426 dvss.n425 0.479667
R906 dvss.n427 dvss.n420 0.479667
R907 dvss.n452 dvss 0.472936
R908 dvss.n439 dvss.n318 0.466883
R909 dvss.n423 dvss.n421 0.451542
R910 dvss.n425 dvss.n424 0.451542
R911 dvss.n422 dvss.n420 0.451542
R912 dvss.n327 dvss.n326 0.440717
R913 dvss.n326 dvss.n325 0.440717
R914 dvss.n383 dvss.n350 0.440717
R915 dvss.n380 dvss.n350 0.440717
R916 dvss.n352 dvss.n351 0.440717
R917 dvss.n353 dvss.n352 0.440717
R918 dvss.n387 dvss.n346 0.440717
R919 dvss.n384 dvss.n346 0.440717
R920 dvss.n348 dvss.n347 0.440717
R921 dvss.n349 dvss.n348 0.440717
R922 dvss.n391 dvss.n342 0.440717
R923 dvss.n388 dvss.n342 0.440717
R924 dvss.n344 dvss.n343 0.440717
R925 dvss.n345 dvss.n344 0.440717
R926 dvss.n341 dvss.n337 0.440717
R927 dvss.n392 dvss.n341 0.440717
R928 dvss.n395 dvss.n339 0.440717
R929 dvss.n340 dvss.n339 0.440717
R930 dvss.n412 dvss.n328 0.440717
R931 dvss.n415 dvss.n328 0.440717
R932 dvss.n331 dvss.n330 0.440717
R933 dvss.n330 dvss.n329 0.440717
R934 dvss.n416 dvss.n324 0.440717
R935 dvss.n419 dvss.n324 0.440717
R936 dvss.n366 dvss.n365 0.440717
R937 dvss.n367 dvss.n366 0.440717
R938 dvss.n369 dvss.n368 0.440717
R939 dvss.n370 dvss.n369 0.440717
R940 dvss.n443 dvss.n442 0.40902
R941 dvss.n448 dvss.n443 0.40902
R942 dvss.n28 dvss.n26 0.38259
R943 dvss.n473 dvss.n454 0.379594
R944 dvss.n496 dvss.n478 0.379594
R945 dvss.n561 dvss.n560 0.379594
R946 dvss.n575 dvss.n2 0.379594
R947 dvss.n451 dvss.n450 0.377433
R948 dvss.n450 dvss.n449 0.377433
R949 dvss.n519 dvss.n515 0.366214
R950 dvss.n359 dvss.n358 0.359196
R951 dvss.n379 dvss.n354 0.359196
R952 dvss.n361 dvss.n354 0.359196
R953 dvss.n397 dvss.n396 0.359196
R954 dvss.n411 dvss.n332 0.359196
R955 dvss.n406 dvss.n334 0.359196
R956 dvss.n403 dvss.n334 0.359196
R957 dvss.n336 dvss.n335 0.359196
R958 dvss.n402 dvss.n336 0.359196
R959 dvss.n398 dvss.n338 0.359196
R960 dvss.n401 dvss.n338 0.359196
R961 dvss.n408 dvss.n407 0.359196
R962 dvss.n407 dvss.n333 0.359196
R963 dvss.n371 dvss.n364 0.359196
R964 dvss.n374 dvss.n364 0.359196
R965 dvss.n363 dvss.n357 0.359196
R966 dvss.n375 dvss.n363 0.359196
R967 dvss.n378 dvss.n356 0.359196
R968 dvss.n362 dvss.n356 0.359196
R969 dvss.n381 dvss.n353 0.351043
R970 dvss.n381 dvss.n380 0.351043
R971 dvss.n382 dvss.n351 0.351043
R972 dvss.n383 dvss.n382 0.351043
R973 dvss.n385 dvss.n349 0.351043
R974 dvss.n385 dvss.n384 0.351043
R975 dvss.n386 dvss.n347 0.351043
R976 dvss.n387 dvss.n386 0.351043
R977 dvss.n389 dvss.n345 0.351043
R978 dvss.n389 dvss.n388 0.351043
R979 dvss.n390 dvss.n343 0.351043
R980 dvss.n391 dvss.n390 0.351043
R981 dvss.n393 dvss.n340 0.351043
R982 dvss.n393 dvss.n392 0.351043
R983 dvss.n395 dvss.n394 0.351043
R984 dvss.n394 dvss.n337 0.351043
R985 dvss.n399 dvss.n398 0.351043
R986 dvss.n409 dvss.n408 0.351043
R987 dvss.n400 dvss.n396 0.351043
R988 dvss.n401 dvss.n400 0.351043
R989 dvss.n410 dvss.n333 0.351043
R990 dvss.n411 dvss.n410 0.351043
R991 dvss.n413 dvss.n331 0.351043
R992 dvss.n413 dvss.n412 0.351043
R993 dvss.n414 dvss.n329 0.351043
R994 dvss.n415 dvss.n414 0.351043
R995 dvss.n417 dvss.n327 0.351043
R996 dvss.n417 dvss.n416 0.351043
R997 dvss.n418 dvss.n325 0.351043
R998 dvss.n419 dvss.n418 0.351043
R999 dvss.n365 dvss.n323 0.351043
R1000 dvss.n367 dvss.n322 0.351043
R1001 dvss.n368 dvss.n321 0.351043
R1002 dvss.n370 dvss.n320 0.351043
R1003 dvss.n358 dvss.n355 0.351043
R1004 dvss.n379 dvss.n355 0.351043
R1005 dvss.n372 dvss.n371 0.351043
R1006 dvss.n361 dvss.n360 0.351043
R1007 dvss.n374 dvss.n373 0.351043
R1008 dvss.n475 dvss.n474 0.332643
R1009 dvss.n498 dvss.n497 0.332643
R1010 dvss.n500 dvss.n14 0.332643
R1011 dvss.n577 dvss.n576 0.332643
R1012 dvss.n441 dvss.n439 0.292684
R1013 dvss.n432 dvss.n323 0.288543
R1014 dvss.n434 dvss.n322 0.288543
R1015 dvss.n435 dvss.n321 0.288543
R1016 dvss.n437 dvss.n320 0.288543
R1017 dvss.n372 dvss.n319 0.288543
R1018 dvss.n373 dvss.n319 0.288543
R1019 dvss.n506 dvss.n505 0.2505
R1020 dvss.n475 dvss 0.242464
R1021 dvss.n498 dvss 0.242464
R1022 dvss.n500 dvss 0.242464
R1023 dvss dvss.n577 0.242464
R1024 dvss.n476 dvss.n475 0.224161
R1025 dvss.n499 dvss.n498 0.224161
R1026 dvss.n501 dvss.n500 0.224161
R1027 dvss.n577 dvss.n0 0.224161
R1028 dvss.n313 dvss.n56 0.217883
R1029 dvss.n441 dvss.n440 0.179826
R1030 dvss.n430 dvss.n428 0.1755
R1031 dvss.n432 dvss.n431 0.120065
R1032 dvss.n440 dvss 0.108642
R1033 dvss.n504 dvss.n476 0.106137
R1034 dvss.n503 dvss.n499 0.106137
R1035 dvss.n502 dvss.n501 0.106137
R1036 dvss.n452 dvss 0.038087
R1037 dvss.n508 dvss.n507 0.0357273
R1038 dvss.n507 dvss.n441 0.0153492
R1039 dvss.n505 dvss 0.0142289
R1040 dvss.n438 dvss.n319 0.00857584
R1041 dvss.n506 dvss.n452 0.000674014
R1042 multiplexer_0.trans_gate_m_31.ena_b multiplexer_0.vtrip_1.t9 97.2843
R1043 multiplexer_0.trans_gate_m_19.ena multiplexer_0.vtrip_1.t2 97.2843
R1044 multiplexer_0.trans_gate_m_31.ena_b multiplexer_0.trans_gate_m_19.ena 19.486
R1045 multiplexer_0.trans_gate_m_31.ena_b multiplexer_0.vtrip_1.t6 18.5516
R1046 multiplexer_0.trans_gate_m_19.ena multiplexer_0.vtrip_1.t4 18.1873
R1047 level_shifter_1.out multiplexer_0.trans_gate_m_31.ena_b 17.2675
R1048 multiplexer_0.vtrip_1.n0 multiplexer_0.vtrip_1.t5 16.8731
R1049 multiplexer_0.trans_gate_m_19.ena multiplexer_0.vtrip_1.t1 16.8731
R1050 multiplexer_0.trans_gate_m_31.ena_b multiplexer_0.vtrip_1.t7 16.8731
R1051 multiplexer_0.vtrip_1.n0 multiplexer_0.vtrip_1.t8 16.5088
R1052 multiplexer_0.trans_gate_m_19.ena multiplexer_0.vtrip_1.t3 16.5088
R1053 multiplexer_0.trans_gate_m_31.ena_b multiplexer_0.vtrip_1.t0 16.5088
R1054 multiplexer_0.trans_gate_m_19.ena multiplexer_0.vtrip_1.n0 14.3239
R1055 multiplexer_0.trans_gate_m_29.in.t3 multiplexer_0.trans_gate_m_29.in.t4 228.216
R1056 multiplexer_0.trans_gate_m_29.in.t3 multiplexer_0.trans_gate_m_29.in.t2 228.216
R1057 multiplexer_0.trans_gate_m_29.in.t3 multiplexer_0.trans_gate_m_29.in.t0 228.216
R1058 multiplexer_0.trans_gate_m_29.in.t3 multiplexer_0.trans_gate_m_29.in.t1 93.7584
R1059 multiplexer_0.trans_gate_m_31.out.t0 multiplexer_0.trans_gate_m_31.out.t4 228.216
R1060 multiplexer_0.trans_gate_m_31.out.t0 multiplexer_0.trans_gate_m_31.out.t3 228.216
R1061 multiplexer_0.trans_gate_m_31.out.t0 multiplexer_0.trans_gate_m_31.out.t1 228.216
R1062 multiplexer_0.trans_gate_m_31.out.t0 multiplexer_0.trans_gate_m_31.out.t2 93.748
R1063 avss.n734 avss.n113 52837.8
R1064 avss.n734 avss.n114 52837.8
R1065 avss.n735 avss.n114 52837.8
R1066 avss.n735 avss.n113 52837.8
R1067 avss.n485 avss.n137 10442.2
R1068 avss.n612 avss.n249 6744.4
R1069 avss.n418 avss.n253 6744.4
R1070 avss.n612 avss.n253 6744.4
R1071 avss.n377 avss.n356 6744.4
R1072 avss.n418 avss.n377 6744.4
R1073 avss.n571 avss.n356 6744.4
R1074 avss.n571 avss.n317 6744.4
R1075 avss.n636 avss.n635 6328.99
R1076 avss.n487 avss.n214 6328.99
R1077 avss.n636 avss.n214 6328.99
R1078 avss.n647 avss.n168 6227.45
R1079 avss.n272 avss.n239 6216.37
R1080 avss.n623 avss.n235 6216.37
R1081 avss.n623 avss.n239 6216.37
R1082 avss.n557 avss.n429 6216.37
R1083 avss.n429 avss.n235 6216.37
R1084 avss.n557 avss.n431 6216.37
R1085 avss.n489 avss.n431 6216.37
R1086 avss.n656 avss.n137 6184.38
R1087 avss.n488 avss.n486 4558.19
R1088 avss.n485 avss.n484 3690.48
R1089 avss.n488 avss.n487 3618.39
R1090 avss.n657 avss.n656 3386.05
R1091 avss.n489 avss.n488 3228.89
R1092 avss.n729 avss.n118 3052.71
R1093 avss.n728 avss.n118 3052.71
R1094 avss.n728 avss.n117 3052.71
R1095 avss.n729 avss.n117 3052.71
R1096 avss.n162 avss.n137 2992.39
R1097 avss.n158 avss.n157 2723.4
R1098 avss.n157 avss.n134 2723.4
R1099 avss.n712 avss.n141 2723.4
R1100 avss.n693 avss.n141 2723.4
R1101 avss.n153 avss.n151 2723.4
R1102 avss.n151 avss.n135 2723.4
R1103 avss.n154 avss.n140 2723.4
R1104 avss.n695 avss.n154 2723.4
R1105 avss.n674 avss.n159 2723.4
R1106 avss.n674 avss.n136 2723.4
R1107 avss.n669 avss.n139 2723.4
R1108 avss.n687 avss.n669 2723.4
R1109 avss.n160 avss.n133 2723.4
R1110 avss.n714 avss.n133 2723.4
R1111 avss.n659 avss.n138 2723.4
R1112 avss.n668 avss.n659 2723.4
R1113 avss.n486 avss.n485 2564.43
R1114 avss.t189 avss.n502 2496.57
R1115 avss.t189 avss.n503 2496.57
R1116 avss.n430 avss.t161 2496.57
R1117 avss.n570 avss.t161 2496.57
R1118 avss.t168 avss.n572 2496.57
R1119 avss.t168 avss.n318 2496.57
R1120 avss.n483 avss.t176 2496.57
R1121 avss.n476 avss.t176 2496.57
R1122 avss.n195 avss.t214 2496.57
R1123 avss.n201 avss.t214 2496.57
R1124 avss.t188 avss.n544 2496.57
R1125 avss.t188 avss.n545 2496.57
R1126 avss.n428 avss.t162 2496.57
R1127 avss.n376 avss.t162 2496.57
R1128 avss.t62 avss.n398 2496.57
R1129 avss.t62 avss.n319 2496.57
R1130 avss.t186 avss.n234 2496.57
R1131 avss.t186 avss.n624 2496.57
R1132 avss.n622 avss.t167 2496.57
R1133 avss.n252 avss.t167 2496.57
R1134 avss.t247 avss.n408 2496.57
R1135 avss.t247 avss.n320 2496.57
R1136 avss.n633 avss.t108 2496.57
R1137 avss.n238 avss.t108 2496.57
R1138 avss.t16 avss.n248 2496.57
R1139 avss.t16 avss.n613 2496.57
R1140 avss.n611 avss.t128 2496.57
R1141 avss.n323 avss.t128 2496.57
R1142 avss.t156 avss.n513 2496.57
R1143 avss.t156 avss.n514 2496.57
R1144 avss.t219 avss.n373 2496.57
R1145 avss.t219 avss.n419 2496.57
R1146 avss.n417 avss.t20 2496.57
R1147 avss.t20 avss.n324 2496.57
R1148 avss.n500 avss.t99 2496.57
R1149 avss.n556 avss.t99 2496.57
R1150 avss.t59 avss.n558 2496.57
R1151 avss.t59 avss.n559 2496.57
R1152 avss.t147 avss.n388 2496.57
R1153 avss.t147 avss.n325 2496.57
R1154 avss.t107 avss.n440 2496.57
R1155 avss.t107 avss.n490 2496.57
R1156 avss.t56 avss.n441 2496.57
R1157 avss.t56 avss.n450 2496.57
R1158 avss.n329 avss.t130 2496.57
R1159 avss.n583 avss.t130 2496.57
R1160 avss.n582 avss.n326 2394.09
R1161 avss.n582 avss.n327 2394.09
R1162 avss.n330 avss.n327 2394.09
R1163 avss.n330 avss.n326 2394.09
R1164 avss.n451 avss.n449 2394.09
R1165 avss.n452 avss.n449 2394.09
R1166 avss.n452 avss.n447 2394.09
R1167 avss.n451 avss.n447 2394.09
R1168 avss.n491 avss.n439 2394.09
R1169 avss.n492 avss.n439 2394.09
R1170 avss.n492 avss.n437 2394.09
R1171 avss.n491 avss.n437 2394.09
R1172 avss.n389 avss.n387 2394.09
R1173 avss.n390 avss.n387 2394.09
R1174 avss.n390 avss.n385 2394.09
R1175 avss.n389 avss.n385 2394.09
R1176 avss.n560 avss.n364 2394.09
R1177 avss.n561 avss.n364 2394.09
R1178 avss.n561 avss.n362 2394.09
R1179 avss.n560 avss.n362 2394.09
R1180 avss.n555 avss.n432 2394.09
R1181 avss.n555 avss.n433 2394.09
R1182 avss.n435 avss.n433 2394.09
R1183 avss.n435 avss.n432 2394.09
R1184 avss.n381 avss.n378 2394.09
R1185 avss.n381 avss.n379 2394.09
R1186 avss.n416 avss.n379 2394.09
R1187 avss.n416 avss.n378 2394.09
R1188 avss.n420 avss.n372 2394.09
R1189 avss.n421 avss.n372 2394.09
R1190 avss.n421 avss.n370 2394.09
R1191 avss.n420 avss.n370 2394.09
R1192 avss.n515 avss.n512 2394.09
R1193 avss.n516 avss.n512 2394.09
R1194 avss.n516 avss.n510 2394.09
R1195 avss.n515 avss.n510 2394.09
R1196 avss.n322 avss.n254 2394.09
R1197 avss.n322 avss.n255 2394.09
R1198 avss.n610 avss.n255 2394.09
R1199 avss.n610 avss.n254 2394.09
R1200 avss.n614 avss.n247 2394.09
R1201 avss.n615 avss.n247 2394.09
R1202 avss.n615 avss.n245 2394.09
R1203 avss.n614 avss.n245 2394.09
R1204 avss.n237 avss.n226 2394.09
R1205 avss.n237 avss.n227 2394.09
R1206 avss.n632 avss.n227 2394.09
R1207 avss.n632 avss.n226 2394.09
R1208 avss.n596 avss.n316 2394.09
R1209 avss.n595 avss.n316 2394.09
R1210 avss.n595 avss.n259 2394.09
R1211 avss.n596 avss.n259 2394.09
R1212 avss.n308 avss.n269 2394.09
R1213 avss.n308 avss.n270 2394.09
R1214 avss.n303 avss.n270 2394.09
R1215 avss.n303 avss.n269 2394.09
R1216 avss.n287 avss.n280 2394.09
R1217 avss.n287 avss.n281 2394.09
R1218 avss.n283 avss.n281 2394.09
R1219 avss.n283 avss.n280 2394.09
R1220 avss.n409 avss.n407 2394.09
R1221 avss.n410 avss.n407 2394.09
R1222 avss.n410 avss.n405 2394.09
R1223 avss.n409 avss.n405 2394.09
R1224 avss.n251 avss.n240 2394.09
R1225 avss.n251 avss.n241 2394.09
R1226 avss.n621 avss.n241 2394.09
R1227 avss.n621 avss.n240 2394.09
R1228 avss.n625 avss.n233 2394.09
R1229 avss.n626 avss.n233 2394.09
R1230 avss.n626 avss.n231 2394.09
R1231 avss.n625 avss.n231 2394.09
R1232 avss.n399 avss.n397 2394.09
R1233 avss.n400 avss.n397 2394.09
R1234 avss.n400 avss.n395 2394.09
R1235 avss.n399 avss.n395 2394.09
R1236 avss.n375 avss.n365 2394.09
R1237 avss.n375 avss.n366 2394.09
R1238 avss.n427 avss.n366 2394.09
R1239 avss.n427 avss.n365 2394.09
R1240 avss.n546 avss.n524 2394.09
R1241 avss.n547 avss.n524 2394.09
R1242 avss.n547 avss.n522 2394.09
R1243 avss.n546 avss.n522 2394.09
R1244 avss.n200 avss.n192 2394.09
R1245 avss.n200 avss.n193 2394.09
R1246 avss.n196 avss.n193 2394.09
R1247 avss.n196 avss.n192 2394.09
R1248 avss.n477 avss.n473 2394.09
R1249 avss.n477 avss.n474 2394.09
R1250 avss.n482 avss.n474 2394.09
R1251 avss.n482 avss.n473 2394.09
R1252 avss.n573 avss.n355 2394.09
R1253 avss.n574 avss.n355 2394.09
R1254 avss.n574 avss.n353 2394.09
R1255 avss.n573 avss.n353 2394.09
R1256 avss.n569 avss.n357 2394.09
R1257 avss.n569 avss.n358 2394.09
R1258 avss.n360 avss.n358 2394.09
R1259 avss.n360 avss.n357 2394.09
R1260 avss.n504 avss.n499 2394.09
R1261 avss.n505 avss.n499 2394.09
R1262 avss.n505 avss.n497 2394.09
R1263 avss.n504 avss.n497 2394.09
R1264 avss.n212 avss.n203 2394.09
R1265 avss.n212 avss.n204 2394.09
R1266 avss.n207 avss.n204 2394.09
R1267 avss.n207 avss.n203 2394.09
R1268 avss.n649 avss.n163 2394.09
R1269 avss.n649 avss.n164 2394.09
R1270 avss.n653 avss.n164 2394.09
R1271 avss.n653 avss.n163 2394.09
R1272 avss.n223 avss.n216 2394.09
R1273 avss.n223 avss.n217 2394.09
R1274 avss.n219 avss.n217 2394.09
R1275 avss.n219 avss.n216 2394.09
R1276 avss.n190 avss.n188 2394.09
R1277 avss.n638 avss.n190 2394.09
R1278 avss.n639 avss.n638 2394.09
R1279 avss.n639 avss.n188 2394.09
R1280 avss.n503 avss.n431 2027.45
R1281 avss.n431 avss.n430 2027.45
R1282 avss.n545 avss.n429 2027.45
R1283 avss.n429 avss.n428 2027.45
R1284 avss.n624 avss.n623 2027.45
R1285 avss.n623 avss.n622 2027.45
R1286 avss.n239 avss.n238 2027.45
R1287 avss.n248 avss.n239 2027.45
R1288 avss.n514 avss.n235 2027.45
R1289 avss.n373 avss.n235 2027.45
R1290 avss.n557 avss.n556 2027.45
R1291 avss.n558 avss.n557 2027.45
R1292 avss.n490 avss.n489 2027.45
R1293 avss.n489 avss.n441 2027.45
R1294 avss.n484 avss.n162 2007.05
R1295 avss.n655 avss.n162 1963.94
R1296 avss.n571 avss.n570 1908.82
R1297 avss.n572 avss.n571 1908.82
R1298 avss.n377 avss.n376 1908.82
R1299 avss.n398 avss.n377 1908.82
R1300 avss.n253 avss.n252 1908.82
R1301 avss.n408 avss.n253 1908.82
R1302 avss.n613 avss.n612 1908.82
R1303 avss.n612 avss.n611 1908.82
R1304 avss.n419 avss.n418 1908.82
R1305 avss.n418 avss.n417 1908.82
R1306 avss.n559 avss.n356 1908.82
R1307 avss.n388 avss.n356 1908.82
R1308 avss.n450 avss.n317 1908.82
R1309 avss.n329 avss.n317 1908.82
R1310 avss.n489 avss.n317 1784.13
R1311 avss.n311 avss.n263 1552.82
R1312 avss.n603 avss.n263 1552.82
R1313 avss.n600 avss.n265 1552.82
R1314 avss.n601 avss.n600 1552.82
R1315 avss.n295 avss.n279 1552.82
R1316 avss.n295 avss.n273 1552.82
R1317 avss.n292 avss.n274 1552.82
R1318 avss.n300 avss.n274 1552.82
R1319 avss.n341 avss.n338 1552.82
R1320 avss.n338 avss.n337 1552.82
R1321 avss.n347 avss.n343 1552.82
R1322 avss.n347 avss.n344 1552.82
R1323 avss.n462 avss.n459 1552.82
R1324 avss.n459 avss.n442 1552.82
R1325 avss.n465 avss.n443 1552.82
R1326 avss.n471 avss.n443 1552.82
R1327 avss.n542 avss.n525 1552.82
R1328 avss.n531 avss.n525 1552.82
R1329 avss.n536 avss.n191 1552.82
R1330 avss.n646 avss.n173 1552.82
R1331 avss.n646 avss.n174 1552.82
R1332 avss.n181 avss.n166 1552.82
R1333 avss.n590 avss.n584 1552.82
R1334 avss.n586 avss.n584 1552.82
R1335 avss.n587 avss.n586 1552.82
R1336 avss.n590 avss.n587 1552.82
R1337 avss.n689 avss.n688 1524.71
R1338 avss.n688 avss.n142 1524.71
R1339 avss.n698 avss.n696 1524.71
R1340 avss.n698 avss.n697 1524.71
R1341 avss.n683 avss.n670 1524.71
R1342 avss.n683 avss.n682 1524.71
R1343 avss.n664 avss.n660 1524.71
R1344 avss.n664 avss.n132 1524.71
R1345 avss.n592 avss.n317 1481.39
R1346 avss.n476 avss.n169 1380.39
R1347 avss.n202 avss.n201 1380.39
R1348 avss.n733 avss.n112 1306.82
R1349 avss.n733 avss.n732 1306.74
R1350 avss.n195 avss.n170 1267.16
R1351 avss.n487 avss.n440 1266.54
R1352 avss.n655 avss.n161 1248.77
R1353 avss.n544 avss.n543 1218.63
R1354 avss.n689 avss.n158 1198.69
R1355 avss.n712 avss.n142 1198.69
R1356 avss.n142 avss.n134 1198.69
R1357 avss.n693 avss.n689 1198.69
R1358 avss.n696 avss.n153 1198.69
R1359 avss.n697 avss.n140 1198.69
R1360 avss.n697 avss.n135 1198.69
R1361 avss.n696 avss.n695 1198.69
R1362 avss.n670 avss.n159 1198.69
R1363 avss.n682 avss.n139 1198.69
R1364 avss.n682 avss.n136 1198.69
R1365 avss.n687 avss.n670 1198.69
R1366 avss.n660 avss.n160 1198.69
R1367 avss.n138 avss.n132 1198.69
R1368 avss.n714 avss.n132 1198.69
R1369 avss.n668 avss.n660 1198.69
R1370 avss.n656 avss.n655 1183.26
R1371 avss.n647 avss.n166 957.487
R1372 avss.n636 avss.n191 929.78
R1373 avss.n486 avss.n168 881.452
R1374 avss.t23 avss.n167 839.736
R1375 avss.t23 avss.n637 839.736
R1376 avss.n206 avss.t24 839.736
R1377 avss.n213 avss.t24 839.736
R1378 avss.n736 avss.n112 815.148
R1379 avss.n311 avss.n268 799.588
R1380 avss.n268 avss.n265 799.588
R1381 avss.n601 avss.n262 799.588
R1382 avss.n603 avss.n262 799.588
R1383 avss.n293 avss.n279 799.588
R1384 avss.n293 avss.n292 799.588
R1385 avss.n300 avss.n275 799.588
R1386 avss.n275 avss.n273 799.588
R1387 avss.n341 avss.n334 799.588
R1388 avss.n343 avss.n334 799.588
R1389 avss.n344 avss.n335 799.588
R1390 avss.n337 avss.n335 799.588
R1391 avss.n466 avss.n462 799.588
R1392 avss.n466 avss.n465 799.588
R1393 avss.n471 avss.n444 799.588
R1394 avss.n444 avss.n442 799.588
R1395 avss.n542 avss.n526 799.588
R1396 avss.n531 avss.n530 799.588
R1397 avss.n530 avss.n191 799.588
R1398 avss.n538 avss.n526 799.588
R1399 avss.n173 avss.n172 799.588
R1400 avss.n180 avss.n174 799.588
R1401 avss.n183 avss.n180 799.588
R1402 avss.n172 avss.n166 799.588
R1403 avss.n268 avss.n267 753.236
R1404 avss.n267 avss.n262 753.236
R1405 avss.n294 avss.n293 753.236
R1406 avss.n294 avss.n275 753.236
R1407 avss.n348 avss.n334 753.236
R1408 avss.n348 avss.n335 753.236
R1409 avss.n467 avss.n466 753.236
R1410 avss.n467 avss.n444 753.236
R1411 avss.n530 avss.n529 753.236
R1412 avss.n529 avss.n526 753.236
R1413 avss.n172 avss.n171 753.236
R1414 avss.n180 avss.n171 753.236
R1415 avss.t131 avss.n336 720.404
R1416 avss.n464 avss.t185 720.404
R1417 avss.n489 avss.n472 709.321
R1418 avss.t129 avss.n170 700.981
R1419 avss.n543 avss.t13 700.981
R1420 avss.n206 avss.n168 680.133
R1421 avss.n637 avss.n636 672.878
R1422 avss.n214 avss.n213 672.878
R1423 avss.n732 avss.n731 663.183
R1424 avss.n647 avss.n169 647.059
R1425 avss.n654 avss.t227 632.672
R1426 avss.n648 avss.t227 632.672
R1427 avss.n636 avss.n202 620.098
R1428 avss.n342 avss.n317 609.572
R1429 avss.n647 avss.n167 554.909
R1430 avss.n538 avss.n537 550.293
R1431 avss.n183 avss.n182 550.293
R1432 avss.n648 avss.n647 513.789
R1433 avss.n502 avss.n501 512.255
R1434 avss.n592 avss.n318 512.255
R1435 avss.n484 avss.n483 512.255
R1436 avss.n592 avss.n319 512.255
R1437 avss.n234 avss.n215 512.255
R1438 avss.n592 avss.n320 512.255
R1439 avss.n634 avss.n633 512.255
R1440 avss.n592 avss.n323 512.255
R1441 avss.n513 avss.n215 512.255
R1442 avss.n592 avss.n324 512.255
R1443 avss.n501 avss.n500 512.255
R1444 avss.n592 avss.n325 512.255
R1445 avss.n592 avss.n583 512.255
R1446 avss.n636 avss.n215 500.577
R1447 avss.n501 avss.n214 500.577
R1448 avss.n658 avss.n657 447.11
R1449 avss.t187 avss.n225 426.997
R1450 avss.n288 avss.t187 426.997
R1451 avss.n302 avss.t123 426.997
R1452 avss.n309 avss.t123 426.997
R1453 avss.t150 avss.n264 426.997
R1454 avss.t150 avss.n593 426.997
R1455 avss.t1 avss 380.286
R1456 avss.t2 avss 380.286
R1457 avss.t0 avss 380.286
R1458 avss.t153 avss.n161 319.26
R1459 avss.n224 avss.t153 319.26
R1460 avss avss.t1 296.784
R1461 avss.t2 avss 296.784
R1462 avss avss.t0 296.784
R1463 avss.n349 avss.n348 292.5
R1464 avss.n348 avss.t131 292.5
R1465 avss.n344 avss.n331 292.5
R1466 avss.n344 avss.n336 292.5
R1467 avss.n337 avss.n332 292.5
R1468 avss.n337 avss.n336 292.5
R1469 avss.n339 avss.n338 292.5
R1470 avss.t131 avss.n338 292.5
R1471 avss.n341 avss.n340 292.5
R1472 avss.n342 avss.n341 292.5
R1473 avss.n345 avss.n343 292.5
R1474 avss.n343 avss.n342 292.5
R1475 avss.n347 avss.n346 292.5
R1476 avss.t131 avss.n347 292.5
R1477 avss.n468 avss.n467 292.5
R1478 avss.n467 avss.t185 292.5
R1479 avss.n471 avss.n470 292.5
R1480 avss.n472 avss.n471 292.5
R1481 avss.n457 avss.n442 292.5
R1482 avss.n472 avss.n442 292.5
R1483 avss.n460 avss.n459 292.5
R1484 avss.n459 avss.t185 292.5
R1485 avss.n462 avss.n461 292.5
R1486 avss.n464 avss.n462 292.5
R1487 avss.n465 avss.n463 292.5
R1488 avss.n465 avss.n464 292.5
R1489 avss.n445 avss.n443 292.5
R1490 avss.n443 avss.t185 292.5
R1491 avss.n539 avss.n538 292.5
R1492 avss.n536 avss.n535 292.5
R1493 avss.n534 avss.n191 292.5
R1494 avss.n178 avss.n166 292.5
R1495 avss.n181 avss.n179 292.5
R1496 avss.n184 avss.n183 292.5
R1497 avss.n176 avss.n171 292.5
R1498 avss.t129 avss.n171 292.5
R1499 avss.n644 avss.n174 292.5
R1500 avss.n174 avss.n170 292.5
R1501 avss.n175 avss.n173 292.5
R1502 avss.n173 avss.n169 292.5
R1503 avss.n646 avss.n645 292.5
R1504 avss.t129 avss.n646 292.5
R1505 avss.n529 avss.n528 292.5
R1506 avss.n529 avss.t13 292.5
R1507 avss.n542 avss.n541 292.5
R1508 avss.n543 avss.n542 292.5
R1509 avss.n532 avss.n531 292.5
R1510 avss.n531 avss.n202 292.5
R1511 avss.n527 avss.n525 292.5
R1512 avss.n525 avss.t13 292.5
R1513 avss.n294 avss.n277 292.5
R1514 avss.t98 avss.n294 292.5
R1515 avss.n300 avss.n299 292.5
R1516 avss.n301 avss.n300 292.5
R1517 avss.n297 avss.n273 292.5
R1518 avss.n301 avss.n273 292.5
R1519 avss.n296 avss.n295 292.5
R1520 avss.n295 avss.t98 292.5
R1521 avss.n279 avss.n278 292.5
R1522 avss.n289 avss.n279 292.5
R1523 avss.n292 avss.n291 292.5
R1524 avss.n292 avss.n289 292.5
R1525 avss.n276 avss.n274 292.5
R1526 avss.t98 avss.n274 292.5
R1527 avss.n267 avss.n260 292.5
R1528 avss.n267 avss.t95 292.5
R1529 avss.n601 avss.n258 292.5
R1530 avss.n602 avss.n601 292.5
R1531 avss.n604 avss.n603 292.5
R1532 avss.n603 avss.n602 292.5
R1533 avss.n266 avss.n263 292.5
R1534 avss.t95 avss.n263 292.5
R1535 avss.n312 avss.n311 292.5
R1536 avss.n311 avss.n310 292.5
R1537 avss.n314 avss.n265 292.5
R1538 avss.n310 avss.n265 292.5
R1539 avss.n600 avss.n599 292.5
R1540 avss.n600 avss.t95 292.5
R1541 avss.n590 avss.n589 292.5
R1542 avss.n591 avss.n590 292.5
R1543 avss.n588 avss.n584 292.5
R1544 avss.n584 avss.t100 292.5
R1545 avss.n586 avss.n123 292.5
R1546 avss.n586 avss.n585 292.5
R1547 avss.n587 avss.n122 292.5
R1548 avss.n587 avss.t100 292.5
R1549 avss.n581 avss.n328 278.212
R1550 avss.n354 avss.n352 278.212
R1551 avss.n386 avss.n384 278.212
R1552 avss.n396 avss.n394 278.212
R1553 avss.n382 avss.n380 278.212
R1554 avss.n406 avss.n404 278.212
R1555 avss.n321 avss.n256 278.212
R1556 avss.n597 avss.n315 278.212
R1557 avss.n448 avss.n446 278.212
R1558 avss.n568 avss.n359 278.212
R1559 avss.n363 avss.n361 278.212
R1560 avss.n374 avss.n367 278.212
R1561 avss.n371 avss.n369 278.212
R1562 avss.n250 avss.n242 278.212
R1563 avss.n246 avss.n244 278.212
R1564 avss.n307 avss.n271 278.212
R1565 avss.n478 avss.n475 278.212
R1566 avss.n650 avss.n165 278.212
R1567 avss.n438 avss.n436 278.212
R1568 avss.n498 avss.n496 278.212
R1569 avss.n554 avss.n434 278.212
R1570 avss.n523 avss.n521 278.212
R1571 avss.n511 avss.n509 278.212
R1572 avss.n232 avss.n230 278.212
R1573 avss.n236 avss.n228 278.212
R1574 avss.n286 avss.n282 278.212
R1575 avss.n222 avss.n218 278.212
R1576 avss.n211 avss.n205 278.212
R1577 avss.n199 avss.n194 278.212
R1578 avss.n189 avss.n186 278.212
R1579 avss.n635 avss.n224 255.822
R1580 avss.n713 avss.t6 241.147
R1581 avss.n302 avss.n301 228.715
R1582 avss.t3 avss 226.321
R1583 avss.n289 avss.n288 225.026
R1584 avss.n310 avss.n309 225.026
R1585 avss.n694 avss.n658 220.312
R1586 avss.n581 avss.n580 214.03
R1587 avss.n575 avss.n354 214.03
R1588 avss.n391 avss.n386 214.03
R1589 avss.n401 avss.n396 214.03
R1590 avss.n383 avss.n382 214.03
R1591 avss.n411 avss.n406 214.03
R1592 avss.n321 avss.n257 214.03
R1593 avss.n594 avss.n315 214.03
R1594 avss.n453 avss.n448 214.03
R1595 avss.n568 avss.n567 214.03
R1596 avss.n562 avss.n363 214.03
R1597 avss.n374 avss.n368 214.03
R1598 avss.n422 avss.n371 214.03
R1599 avss.n250 avss.n243 214.03
R1600 avss.n616 avss.n246 214.03
R1601 avss.n307 avss.n306 214.03
R1602 avss.n479 avss.n478 214.03
R1603 avss.n651 avss.n650 214.03
R1604 avss.n493 avss.n438 214.03
R1605 avss.n506 avss.n498 214.03
R1606 avss.n554 avss.n553 214.03
R1607 avss.n548 avss.n523 214.03
R1608 avss.n517 avss.n511 214.03
R1609 avss.n627 avss.n232 214.03
R1610 avss.n236 avss.n229 214.03
R1611 avss.n286 avss.n285 214.03
R1612 avss.n222 avss.n221 214.03
R1613 avss.n211 avss.n210 214.03
R1614 avss.n199 avss.n198 214.03
R1615 avss.n189 avss.n187 214.03
R1616 avss.n579 avss.n328 204.909
R1617 avss.n576 avss.n352 204.909
R1618 avss.n392 avss.n384 204.909
R1619 avss.n402 avss.n394 204.909
R1620 avss.n415 avss.n380 204.909
R1621 avss.n412 avss.n404 204.909
R1622 avss.n609 avss.n256 204.909
R1623 avss.n454 avss.n446 204.909
R1624 avss.n566 avss.n359 204.909
R1625 avss.n563 avss.n361 204.909
R1626 avss.n426 avss.n367 204.909
R1627 avss.n423 avss.n369 204.909
R1628 avss.n620 avss.n242 204.909
R1629 avss.n617 avss.n244 204.909
R1630 avss.n305 avss.n271 204.909
R1631 avss.n481 avss.n475 204.909
R1632 avss.n652 avss.n165 204.909
R1633 avss.n494 avss.n436 204.909
R1634 avss.n507 avss.n496 204.909
R1635 avss.n552 avss.n434 204.909
R1636 avss.n549 avss.n521 204.909
R1637 avss.n518 avss.n509 204.909
R1638 avss.n628 avss.n230 204.909
R1639 avss.n631 avss.n228 204.909
R1640 avss.n284 avss.n282 204.909
R1641 avss.n220 avss.n218 204.909
R1642 avss.n209 avss.n205 204.909
R1643 avss.n197 avss.n194 204.909
R1644 avss.n640 avss.n186 204.909
R1645 avss.n635 avss.n634 190.315
R1646 avss.n602 avss.n264 188.137
R1647 avss.n598 avss.n597 187.107
R1648 avss.n655 avss.n654 183.107
R1649 avss.n691 avss.n144 174.306
R1650 avss.n710 avss.n144 174.306
R1651 avss.n699 avss.n150 174.306
R1652 avss.n700 avss.n699 174.306
R1653 avss.n685 avss.n684 174.306
R1654 avss.n684 avss.n681 174.306
R1655 avss.n666 avss.n665 174.306
R1656 avss.n665 avss.n131 174.306
R1657 avss.n711 avss.n143 170.748
R1658 avss.n692 avss.n143 170.748
R1659 avss.n155 avss.n149 170.748
R1660 avss.n156 avss.n155 170.748
R1661 avss.n673 avss.n671 170.748
R1662 avss.n686 avss.n671 170.748
R1663 avss.n662 avss.n661 170.748
R1664 avss.n667 avss.n662 170.748
R1665 avss.n690 avss.n145 166.988
R1666 avss.n152 avss.n148 166.988
R1667 avss.n675 avss.n672 166.988
R1668 avss.n663 avss.n130 166.988
R1669 avss.n709 avss.n708 166.934
R1670 avss.n702 avss.n701 166.934
R1671 avss.n680 avss.n679 166.934
R1672 avss.n716 avss.n715 166.934
R1673 avss.n537 avss.n536 158.911
R1674 avss.n182 avss.n181 158.911
R1675 avss.t8 avss.n114 145.641
R1676 avss.n120 avss.t3 143.45
R1677 avss avss.t8 142.819
R1678 avss.n711 avss.n710 141.554
R1679 avss.n692 avss.n691 141.554
R1680 avss.n691 avss.n690 141.554
R1681 avss.n710 avss.n709 141.554
R1682 avss.n700 avss.n149 141.554
R1683 avss.n156 avss.n150 141.554
R1684 avss.n152 avss.n150 141.554
R1685 avss.n701 avss.n700 141.554
R1686 avss.n681 avss.n673 141.554
R1687 avss.n686 avss.n685 141.554
R1688 avss.n685 avss.n672 141.554
R1689 avss.n681 avss.n680 141.554
R1690 avss.n666 avss.n663 141.554
R1691 avss.n661 avss.n131 141.554
R1692 avss.n715 avss.n131 141.554
R1693 avss.n667 avss.n666 141.554
R1694 avss.t98 avss.n289 119.891
R1695 avss.n602 avss.t95 119.891
R1696 avss.n301 avss.n272 118.047
R1697 avss.n580 avss.n579 117.334
R1698 avss.n576 avss.n575 117.334
R1699 avss.n392 avss.n391 117.334
R1700 avss.n402 avss.n401 117.334
R1701 avss.n415 avss.n383 117.334
R1702 avss.n412 avss.n411 117.334
R1703 avss.n609 avss.n257 117.334
R1704 avss.n454 avss.n453 117.334
R1705 avss.n567 avss.n566 117.334
R1706 avss.n563 avss.n562 117.334
R1707 avss.n426 avss.n368 117.334
R1708 avss.n423 avss.n422 117.334
R1709 avss.n620 avss.n243 117.334
R1710 avss.n617 avss.n616 117.334
R1711 avss.n306 avss.n305 117.334
R1712 avss.n481 avss.n479 117.334
R1713 avss.n652 avss.n651 117.334
R1714 avss.n494 avss.n493 117.334
R1715 avss.n507 avss.n506 117.334
R1716 avss.n553 avss.n552 117.334
R1717 avss.n549 avss.n548 117.334
R1718 avss.n518 avss.n517 117.334
R1719 avss.n628 avss.n627 117.334
R1720 avss.n631 avss.n229 117.334
R1721 avss.n285 avss.n284 117.334
R1722 avss.n221 avss.n220 117.334
R1723 avss.n210 avss.n209 117.334
R1724 avss.n198 avss.n197 117.334
R1725 avss.n640 avss.n187 117.334
R1726 avss.t131 avss.n317 110.832
R1727 avss.n537 avss.t19 103.657
R1728 avss.n182 avss.t250 103.657
R1729 avss.n310 avss.n249 101.447
R1730 avss.n599 avss.n314 100.894
R1731 avss.n312 avss.n266 100.894
R1732 avss.n340 avss.n339 100.894
R1733 avss.n346 avss.n345 100.894
R1734 avss.n291 avss.n276 100.894
R1735 avss.n296 avss.n278 100.894
R1736 avss.n461 avss.n460 100.894
R1737 avss.n463 avss.n445 100.894
R1738 avss.n532 avss.n527 100.894
R1739 avss.n535 avss.n534 100.894
R1740 avss.n645 avss.n175 100.894
R1741 avss.n179 avss.n178 100.894
R1742 avss.n640 avss.n639 97.5005
R1743 avss.n639 avss.n167 97.5005
R1744 avss.n190 avss.n189 97.5005
R1745 avss.n637 avss.n190 97.5005
R1746 avss.n220 avss.n219 97.5005
R1747 avss.n219 avss.n161 97.5005
R1748 avss.n223 avss.n222 97.5005
R1749 avss.n224 avss.n223 97.5005
R1750 avss.n653 avss.n652 97.5005
R1751 avss.n654 avss.n653 97.5005
R1752 avss.n650 avss.n649 97.5005
R1753 avss.n649 avss.n648 97.5005
R1754 avss.n209 avss.n207 97.5005
R1755 avss.n207 avss.n206 97.5005
R1756 avss.n212 avss.n211 97.5005
R1757 avss.n213 avss.n212 97.5005
R1758 avss.n507 avss.n497 97.5005
R1759 avss.n502 avss.n497 97.5005
R1760 avss.n499 avss.n498 97.5005
R1761 avss.n503 avss.n499 97.5005
R1762 avss.n566 avss.n360 97.5005
R1763 avss.n430 avss.n360 97.5005
R1764 avss.n569 avss.n568 97.5005
R1765 avss.n570 avss.n569 97.5005
R1766 avss.n576 avss.n353 97.5005
R1767 avss.n572 avss.n353 97.5005
R1768 avss.n355 avss.n354 97.5005
R1769 avss.n355 avss.n318 97.5005
R1770 avss.n482 avss.n481 97.5005
R1771 avss.n483 avss.n482 97.5005
R1772 avss.n478 avss.n477 97.5005
R1773 avss.n477 avss.n476 97.5005
R1774 avss.n197 avss.n196 97.5005
R1775 avss.n196 avss.n195 97.5005
R1776 avss.n200 avss.n199 97.5005
R1777 avss.n201 avss.n200 97.5005
R1778 avss.n549 avss.n522 97.5005
R1779 avss.n544 avss.n522 97.5005
R1780 avss.n524 avss.n523 97.5005
R1781 avss.n545 avss.n524 97.5005
R1782 avss.n427 avss.n426 97.5005
R1783 avss.n428 avss.n427 97.5005
R1784 avss.n375 avss.n374 97.5005
R1785 avss.n376 avss.n375 97.5005
R1786 avss.n402 avss.n395 97.5005
R1787 avss.n398 avss.n395 97.5005
R1788 avss.n397 avss.n396 97.5005
R1789 avss.n397 avss.n319 97.5005
R1790 avss.n628 avss.n231 97.5005
R1791 avss.n234 avss.n231 97.5005
R1792 avss.n233 avss.n232 97.5005
R1793 avss.n624 avss.n233 97.5005
R1794 avss.n621 avss.n620 97.5005
R1795 avss.n622 avss.n621 97.5005
R1796 avss.n251 avss.n250 97.5005
R1797 avss.n252 avss.n251 97.5005
R1798 avss.n412 avss.n405 97.5005
R1799 avss.n408 avss.n405 97.5005
R1800 avss.n407 avss.n406 97.5005
R1801 avss.n407 avss.n320 97.5005
R1802 avss.n284 avss.n283 97.5005
R1803 avss.n283 avss.n225 97.5005
R1804 avss.n287 avss.n286 97.5005
R1805 avss.n288 avss.n287 97.5005
R1806 avss.n305 avss.n303 97.5005
R1807 avss.n303 avss.n302 97.5005
R1808 avss.n308 avss.n307 97.5005
R1809 avss.n309 avss.n308 97.5005
R1810 avss.n606 avss.n259 97.5005
R1811 avss.n264 avss.n259 97.5005
R1812 avss.n316 avss.n315 97.5005
R1813 avss.n593 avss.n316 97.5005
R1814 avss.n632 avss.n631 97.5005
R1815 avss.n633 avss.n632 97.5005
R1816 avss.n237 avss.n236 97.5005
R1817 avss.n238 avss.n237 97.5005
R1818 avss.n617 avss.n245 97.5005
R1819 avss.n248 avss.n245 97.5005
R1820 avss.n247 avss.n246 97.5005
R1821 avss.n613 avss.n247 97.5005
R1822 avss.n610 avss.n609 97.5005
R1823 avss.n611 avss.n610 97.5005
R1824 avss.n322 avss.n321 97.5005
R1825 avss.n323 avss.n322 97.5005
R1826 avss.n518 avss.n510 97.5005
R1827 avss.n513 avss.n510 97.5005
R1828 avss.n512 avss.n511 97.5005
R1829 avss.n514 avss.n512 97.5005
R1830 avss.n423 avss.n370 97.5005
R1831 avss.n373 avss.n370 97.5005
R1832 avss.n372 avss.n371 97.5005
R1833 avss.n419 avss.n372 97.5005
R1834 avss.n416 avss.n415 97.5005
R1835 avss.n417 avss.n416 97.5005
R1836 avss.n382 avss.n381 97.5005
R1837 avss.n381 avss.n324 97.5005
R1838 avss.n552 avss.n435 97.5005
R1839 avss.n500 avss.n435 97.5005
R1840 avss.n555 avss.n554 97.5005
R1841 avss.n556 avss.n555 97.5005
R1842 avss.n563 avss.n362 97.5005
R1843 avss.n558 avss.n362 97.5005
R1844 avss.n364 avss.n363 97.5005
R1845 avss.n559 avss.n364 97.5005
R1846 avss.n392 avss.n385 97.5005
R1847 avss.n388 avss.n385 97.5005
R1848 avss.n387 avss.n386 97.5005
R1849 avss.n387 avss.n325 97.5005
R1850 avss.n494 avss.n437 97.5005
R1851 avss.n440 avss.n437 97.5005
R1852 avss.n439 avss.n438 97.5005
R1853 avss.n490 avss.n439 97.5005
R1854 avss.n454 avss.n447 97.5005
R1855 avss.n447 avss.n441 97.5005
R1856 avss.n449 avss.n448 97.5005
R1857 avss.n450 avss.n449 97.5005
R1858 avss.n579 avss.n330 97.5005
R1859 avss.n330 avss.n329 97.5005
R1860 avss.n582 avss.n581 97.5005
R1861 avss.n583 avss.n582 97.5005
R1862 avss.t223 avss.n119 97.3856
R1863 avss.t223 avss.n121 97.3856
R1864 avss.n594 avss.n261 95.7798
R1865 avss.n634 avss.n225 87.6132
R1866 avss.n593 avss.n592 87.6132
R1867 avss.n636 avss.t19 83.1239
R1868 avss.n636 avss.t13 80.8829
R1869 avss.n541 avss.n527 72.1417
R1870 avss.n539 avss.n535 72.1417
R1871 avss.n645 avss.n644 68.4924
R1872 avss.n184 avss.n179 68.4924
R1873 avss.n339 avss.n332 67.468
R1874 avss.n346 avss.n331 67.468
R1875 avss.n299 avss.n276 67.468
R1876 avss.n297 avss.n296 67.468
R1877 avss.n460 avss.n457 67.468
R1878 avss.n470 avss.n445 67.468
R1879 avss.n668 avss.n667 65.0005
R1880 avss.n694 avss.n668 65.0005
R1881 avss.n661 avss.n138 65.0005
R1882 avss.n713 avss.n138 65.0005
R1883 avss.n663 avss.n160 65.0005
R1884 avss.n694 avss.n160 65.0005
R1885 avss.n715 avss.n714 65.0005
R1886 avss.n714 avss.n713 65.0005
R1887 avss.n687 avss.n686 65.0005
R1888 avss.n694 avss.n687 65.0005
R1889 avss.n673 avss.n139 65.0005
R1890 avss.n713 avss.n139 65.0005
R1891 avss.n672 avss.n159 65.0005
R1892 avss.n694 avss.n159 65.0005
R1893 avss.n680 avss.n136 65.0005
R1894 avss.n713 avss.n136 65.0005
R1895 avss.n695 avss.n156 65.0005
R1896 avss.n695 avss.n694 65.0005
R1897 avss.n149 avss.n140 65.0005
R1898 avss.n713 avss.n140 65.0005
R1899 avss.n153 avss.n152 65.0005
R1900 avss.n694 avss.n153 65.0005
R1901 avss.n701 avss.n135 65.0005
R1902 avss.n713 avss.n135 65.0005
R1903 avss.n693 avss.n692 65.0005
R1904 avss.n694 avss.n693 65.0005
R1905 avss.n712 avss.n711 65.0005
R1906 avss.n713 avss.n712 65.0005
R1907 avss.n690 avss.n158 65.0005
R1908 avss.n694 avss.n158 65.0005
R1909 avss.n709 avss.n134 65.0005
R1910 avss.n713 avss.n134 65.0005
R1911 avss.n737 avss.n111 62.759
R1912 avss.n730 avss.n116 61.5669
R1913 avss.n713 avss.n137 59.8963
R1914 avss.n731 avss.n730 59.0984
R1915 avss.n647 avss.t250 55.4161
R1916 avss.n647 avss.t129 53.9221
R1917 avss.n662 avss.n659 53.1823
R1918 avss.n659 avss.t6 53.1823
R1919 avss.n665 avss.n664 53.1823
R1920 avss.n664 avss.t6 53.1823
R1921 avss.n671 avss.n669 53.1823
R1922 avss.n669 avss.t6 53.1823
R1923 avss.n684 avss.n683 53.1823
R1924 avss.n683 avss.t6 53.1823
R1925 avss.n675 avss.n674 53.1823
R1926 avss.n674 avss.t6 53.1823
R1927 avss.n155 avss.n154 53.1823
R1928 avss.n154 avss.t6 53.1823
R1929 avss.n699 avss.n698 53.1823
R1930 avss.n698 avss.t6 53.1823
R1931 avss.n151 avss.n148 53.1823
R1932 avss.n151 avss.t6 53.1823
R1933 avss.n143 avss.n141 53.1823
R1934 avss.n141 avss.t6 53.1823
R1935 avss.n688 avss.n144 53.1823
R1936 avss.n688 avss.t6 53.1823
R1937 avss.n157 avss.n145 53.1823
R1938 avss.n157 avss.t6 53.1823
R1939 avss.n133 avss.n130 53.1823
R1940 avss.n657 avss.n133 53.1823
R1941 avss.n188 avss.n186 53.1823
R1942 avss.t23 avss.n188 53.1823
R1943 avss.n638 avss.n187 53.1823
R1944 avss.n638 avss.t23 53.1823
R1945 avss.n218 avss.n216 53.1823
R1946 avss.n216 avss.t153 53.1823
R1947 avss.n221 avss.n217 53.1823
R1948 avss.n217 avss.t153 53.1823
R1949 avss.n165 avss.n163 53.1823
R1950 avss.n163 avss.t227 53.1823
R1951 avss.n651 avss.n164 53.1823
R1952 avss.n164 avss.t227 53.1823
R1953 avss.n205 avss.n203 53.1823
R1954 avss.n203 avss.t24 53.1823
R1955 avss.n210 avss.n204 53.1823
R1956 avss.n204 avss.t24 53.1823
R1957 avss.n504 avss.n496 53.1823
R1958 avss.t189 avss.n504 53.1823
R1959 avss.n506 avss.n505 53.1823
R1960 avss.n505 avss.t189 53.1823
R1961 avss.n359 avss.n357 53.1823
R1962 avss.n357 avss.t161 53.1823
R1963 avss.n567 avss.n358 53.1823
R1964 avss.n358 avss.t161 53.1823
R1965 avss.n573 avss.n352 53.1823
R1966 avss.t168 avss.n573 53.1823
R1967 avss.n575 avss.n574 53.1823
R1968 avss.n574 avss.t168 53.1823
R1969 avss.n475 avss.n473 53.1823
R1970 avss.n473 avss.t176 53.1823
R1971 avss.n479 avss.n474 53.1823
R1972 avss.n474 avss.t176 53.1823
R1973 avss.n194 avss.n192 53.1823
R1974 avss.n192 avss.t214 53.1823
R1975 avss.n198 avss.n193 53.1823
R1976 avss.n193 avss.t214 53.1823
R1977 avss.n546 avss.n521 53.1823
R1978 avss.t188 avss.n546 53.1823
R1979 avss.n548 avss.n547 53.1823
R1980 avss.n547 avss.t188 53.1823
R1981 avss.n367 avss.n365 53.1823
R1982 avss.n365 avss.t162 53.1823
R1983 avss.n368 avss.n366 53.1823
R1984 avss.n366 avss.t162 53.1823
R1985 avss.n399 avss.n394 53.1823
R1986 avss.t62 avss.n399 53.1823
R1987 avss.n401 avss.n400 53.1823
R1988 avss.n400 avss.t62 53.1823
R1989 avss.n625 avss.n230 53.1823
R1990 avss.t186 avss.n625 53.1823
R1991 avss.n627 avss.n626 53.1823
R1992 avss.n626 avss.t186 53.1823
R1993 avss.n242 avss.n240 53.1823
R1994 avss.n240 avss.t167 53.1823
R1995 avss.n243 avss.n241 53.1823
R1996 avss.n241 avss.t167 53.1823
R1997 avss.n409 avss.n404 53.1823
R1998 avss.t247 avss.n409 53.1823
R1999 avss.n411 avss.n410 53.1823
R2000 avss.n410 avss.t247 53.1823
R2001 avss.n282 avss.n280 53.1823
R2002 avss.n280 avss.t187 53.1823
R2003 avss.n285 avss.n281 53.1823
R2004 avss.n281 avss.t187 53.1823
R2005 avss.n271 avss.n269 53.1823
R2006 avss.n269 avss.t123 53.1823
R2007 avss.n306 avss.n270 53.1823
R2008 avss.n270 avss.t123 53.1823
R2009 avss.n597 avss.n596 53.1823
R2010 avss.n596 avss.t150 53.1823
R2011 avss.n595 avss.n594 53.1823
R2012 avss.t150 avss.n595 53.1823
R2013 avss.n228 avss.n226 53.1823
R2014 avss.n226 avss.t108 53.1823
R2015 avss.n229 avss.n227 53.1823
R2016 avss.n227 avss.t108 53.1823
R2017 avss.n614 avss.n244 53.1823
R2018 avss.t16 avss.n614 53.1823
R2019 avss.n616 avss.n615 53.1823
R2020 avss.n615 avss.t16 53.1823
R2021 avss.n256 avss.n254 53.1823
R2022 avss.n254 avss.t128 53.1823
R2023 avss.n257 avss.n255 53.1823
R2024 avss.n255 avss.t128 53.1823
R2025 avss.n515 avss.n509 53.1823
R2026 avss.t156 avss.n515 53.1823
R2027 avss.n517 avss.n516 53.1823
R2028 avss.n516 avss.t156 53.1823
R2029 avss.n420 avss.n369 53.1823
R2030 avss.t219 avss.n420 53.1823
R2031 avss.n422 avss.n421 53.1823
R2032 avss.n421 avss.t219 53.1823
R2033 avss.n380 avss.n378 53.1823
R2034 avss.n378 avss.t20 53.1823
R2035 avss.n383 avss.n379 53.1823
R2036 avss.n379 avss.t20 53.1823
R2037 avss.n434 avss.n432 53.1823
R2038 avss.n432 avss.t99 53.1823
R2039 avss.n553 avss.n433 53.1823
R2040 avss.n433 avss.t99 53.1823
R2041 avss.n560 avss.n361 53.1823
R2042 avss.t59 avss.n560 53.1823
R2043 avss.n562 avss.n561 53.1823
R2044 avss.n561 avss.t59 53.1823
R2045 avss.n389 avss.n384 53.1823
R2046 avss.t147 avss.n389 53.1823
R2047 avss.n391 avss.n390 53.1823
R2048 avss.n390 avss.t147 53.1823
R2049 avss.n491 avss.n436 53.1823
R2050 avss.t107 avss.n491 53.1823
R2051 avss.n493 avss.n492 53.1823
R2052 avss.n492 avss.t107 53.1823
R2053 avss.n451 avss.n446 53.1823
R2054 avss.t56 avss.n451 53.1823
R2055 avss.n453 avss.n452 53.1823
R2056 avss.n452 avss.t56 53.1823
R2057 avss.n328 avss.n326 53.1823
R2058 avss.n326 avss.t130 53.1823
R2059 avss.n580 avss.n327 53.1823
R2060 avss.n327 avss.t130 53.1823
R2061 avss.n730 avss.n729 53.1823
R2062 avss.n729 avss.t223 53.1823
R2063 avss.n728 avss.n727 53.1823
R2064 avss.t223 avss.n728 53.1823
R2065 avss.n314 avss.n313 51.9534
R2066 avss.n313 avss.n312 51.9534
R2067 avss.n345 avss.n333 51.9534
R2068 avss.n340 avss.n333 51.9534
R2069 avss.n291 avss.n290 51.9534
R2070 avss.n290 avss.n278 51.9534
R2071 avss.n463 avss.n458 51.9534
R2072 avss.n461 avss.n458 51.9534
R2073 avss.n533 avss.n532 51.9534
R2074 avss.n534 avss.n533 51.9534
R2075 avss.n177 avss.n175 51.9534
R2076 avss.n178 avss.n177 51.9534
R2077 avss.n599 avss.n598 50.6259
R2078 avss.n313 avss.n260 48.9417
R2079 avss.n349 avss.n333 48.9417
R2080 avss.n290 avss.n277 48.9417
R2081 avss.n468 avss.n458 48.9417
R2082 avss.n533 avss.n528 48.9417
R2083 avss.n177 avss.n176 48.9417
R2084 avss.n118 avss.n115 48.7505
R2085 avss.n121 avss.n118 48.7505
R2086 avss.n123 avss.n117 48.7505
R2087 avss.n119 avss.n117 48.7505
R2088 avss.n266 avss.n261 43.6169
R2089 avss.n605 avss.n260 42.5417
R2090 avss.n350 avss.n349 42.5417
R2091 avss.n298 avss.n277 42.5417
R2092 avss.n469 avss.n468 42.5417
R2093 avss.n540 avss.n528 42.5417
R2094 avss.n643 avss.n176 42.5417
R2095 avss.n146 avss.t25 41.586
R2096 avss.n147 avss.t169 41.586
R2097 avss.n676 avss.t132 41.586
R2098 avss.n129 avss.t72 41.586
R2099 avss.n146 avss.t222 40.9588
R2100 avss.n147 avss.t69 40.9588
R2101 avss.n676 avss.t7 40.9588
R2102 avss.n129 avss.t240 40.9588
R2103 avss.n731 avss.n115 32.2212
R2104 avss.n589 avss.n122 31.0458
R2105 avss.n541 avss.n540 31.0005
R2106 avss.n540 avss.n539 31.0005
R2107 avss.n725 avss.t224 30.1756
R2108 avss.n589 avss.n588 29.7453
R2109 avss.n591 avss.t100 27.3441
R2110 avss.n585 avss.t100 27.3441
R2111 avss.n644 avss.n643 27.1786
R2112 avss.n643 avss.n184 27.1786
R2113 avss.n115 avss.n111 27.1769
R2114 avss.n350 avss.n331 26.1058
R2115 avss.n350 avss.n332 26.1058
R2116 avss.n299 avss.n298 26.1058
R2117 avss.n298 avss.n297 26.1058
R2118 avss.n470 avss.n469 26.1058
R2119 avss.n469 avss.n457 26.1058
R2120 avss.n585 avss.n119 24.3994
R2121 avss.n121 avss.n120 23.558
R2122 avss.n658 avss.t6 19.4289
R2123 avss.t95 avss.n249 18.4453
R2124 avss.n726 avss.n123 16.7152
R2125 avss.n737 avss.n736 11.7731
R2126 avss.n489 avss.t185 11.0836
R2127 avss.n123 avss.n116 10.9042
R2128 avss.n105 avss.t110 10.7251
R2129 avss.n4 avss.t196 10.6793
R2130 avss.n107 avss.t239 10.5739
R2131 avss.n109 avss.t76 10.5739
R2132 avss.n1 avss.t88 10.5739
R2133 avss.n3 avss.t197 10.5739
R2134 avss.n58 avss.t199 10.5739
R2135 avss.n57 avss.t218 10.5739
R2136 avss.n55 avss.t66 10.5739
R2137 avss.n53 avss.t134 10.5739
R2138 avss.n51 avss.t122 10.5739
R2139 avss.n50 avss.t49 10.5739
R2140 avss.n49 avss.t29 10.5739
R2141 avss.n48 avss.t254 10.5739
R2142 avss.n47 avss.t39 10.5739
R2143 avss.n46 avss.t12 10.5739
R2144 avss.n45 avss.t211 10.5739
R2145 avss.n44 avss.t138 10.5739
R2146 avss.n43 avss.t205 10.5739
R2147 avss.n42 avss.t61 10.5739
R2148 avss.n41 avss.t249 10.5739
R2149 avss.n40 avss.t71 10.5739
R2150 avss.n39 avss.t231 10.5739
R2151 avss.n38 avss.t125 10.5739
R2152 avss.n37 avss.t64 10.5739
R2153 avss.n36 avss.t213 10.5739
R2154 avss.n35 avss.t229 10.5739
R2155 avss.n34 avss.t102 10.5739
R2156 avss.n33 avss.t116 10.5739
R2157 avss.n32 avss.t237 10.5739
R2158 avss.n31 avss.t127 10.5739
R2159 avss.n30 avss.t201 10.5739
R2160 avss.n29 avss.t136 10.5739
R2161 avss.n28 avss.t158 10.5739
R2162 avss.n27 avss.t171 10.5739
R2163 avss.n26 avss.t144 10.5739
R2164 avss.n25 avss.t209 10.5739
R2165 avss.n24 avss.t178 10.5739
R2166 avss.n23 avss.t80 10.5739
R2167 avss.n22 avss.t94 10.5739
R2168 avss.n21 avss.t112 10.5739
R2169 avss.n20 avss.t120 10.5739
R2170 avss.n19 avss.t207 10.5739
R2171 avss.n18 avss.t5 10.5739
R2172 avss.n17 avss.t106 10.5739
R2173 avss.n16 avss.t146 10.5739
R2174 avss.n15 avss.t74 10.5739
R2175 avss.n14 avss.t182 10.5739
R2176 avss.n13 avss.t140 10.5739
R2177 avss.n12 avss.t37 10.5739
R2178 avss.n11 avss.t15 10.5739
R2179 avss.n10 avss.t41 10.5739
R2180 avss.n9 avss.t256 10.5739
R2181 avss.n8 avss.t184 10.5739
R2182 avss.n7 avss.t166 10.5739
R2183 avss.n6 avss.t216 10.5739
R2184 avss.n5 avss.t92 10.5739
R2185 avss.n59 avss.t45 10.5739
R2186 avss.n60 avss.t242 10.5739
R2187 avss.n61 avss.t53 10.5739
R2188 avss.n62 avss.t252 10.5739
R2189 avss.n63 avss.t31 10.5739
R2190 avss.n64 avss.t51 10.5739
R2191 avss.n65 avss.t173 10.5739
R2192 avss.n66 avss.t152 10.5739
R2193 avss.n67 avss.t10 10.5739
R2194 avss.n68 avss.t78 10.5739
R2195 avss.n69 avss.t58 10.5739
R2196 avss.n70 avss.t221 10.5739
R2197 avss.n71 avss.t35 10.5739
R2198 avss.n72 avss.t149 10.5739
R2199 avss.n73 avss.t86 10.5739
R2200 avss.n74 avss.t160 10.5739
R2201 avss.n75 avss.t68 10.5739
R2202 avss.n76 avss.t82 10.5739
R2203 avss.n77 avss.t226 10.5739
R2204 avss.n78 avss.t114 10.5739
R2205 avss.n79 avss.t118 10.5739
R2206 avss.n80 avss.t246 10.5739
R2207 avss.n81 avss.t193 10.5739
R2208 avss.n82 avss.t155 10.5739
R2209 avss.n83 avss.t47 10.5739
R2210 avss.n84 avss.t33 10.5739
R2211 avss.n85 avss.t191 10.5739
R2212 avss.n86 avss.t43 10.5739
R2213 avss.n87 avss.t244 10.5739
R2214 avss.n88 avss.t233 10.5739
R2215 avss.n89 avss.t180 10.5739
R2216 avss.n90 avss.t142 10.5739
R2217 avss.n91 avss.t164 10.5739
R2218 avss.n92 avss.t203 10.5739
R2219 avss.n93 avss.t27 10.5739
R2220 avss.n94 avss.t97 10.5739
R2221 avss.n95 avss.t22 10.5739
R2222 avss.n96 avss.t55 10.5739
R2223 avss.n97 avss.t195 10.5739
R2224 avss.n98 avss.t235 10.5739
R2225 avss.n99 avss.t104 10.5739
R2226 avss.n100 avss.t90 10.5739
R2227 avss.n101 avss.t258 10.5739
R2228 avss.n102 avss.t84 10.5739
R2229 avss.n103 avss.t175 10.5739
R2230 avss.n104 avss.t18 10.5739
R2231 avss.n5 avss.t91 10.5285
R2232 avss.n6 avss.t215 10.5285
R2233 avss.n7 avss.t165 10.5285
R2234 avss.n8 avss.t183 10.5285
R2235 avss.n9 avss.t255 10.5285
R2236 avss.n10 avss.t40 10.5285
R2237 avss.n11 avss.t14 10.5285
R2238 avss.n12 avss.t36 10.5285
R2239 avss.n13 avss.t139 10.5285
R2240 avss.n14 avss.t181 10.5285
R2241 avss.n15 avss.t73 10.5285
R2242 avss.n16 avss.t145 10.5285
R2243 avss.n17 avss.t105 10.5285
R2244 avss.n18 avss.t4 10.5285
R2245 avss.n19 avss.t206 10.5285
R2246 avss.n20 avss.t119 10.5285
R2247 avss.n21 avss.t111 10.5285
R2248 avss.n22 avss.t93 10.5285
R2249 avss.n23 avss.t79 10.5285
R2250 avss.n24 avss.t177 10.5285
R2251 avss.n25 avss.t208 10.5285
R2252 avss.n26 avss.t143 10.5285
R2253 avss.n27 avss.t170 10.5285
R2254 avss.n28 avss.t157 10.5285
R2255 avss.n29 avss.t135 10.5285
R2256 avss.n30 avss.t200 10.5285
R2257 avss.n31 avss.t126 10.5285
R2258 avss.n32 avss.t236 10.5285
R2259 avss.n33 avss.t115 10.5285
R2260 avss.n34 avss.t101 10.5285
R2261 avss.n35 avss.t228 10.5285
R2262 avss.n36 avss.t212 10.5285
R2263 avss.n37 avss.t63 10.5285
R2264 avss.n38 avss.t124 10.5285
R2265 avss.n39 avss.t230 10.5285
R2266 avss.n40 avss.t70 10.5285
R2267 avss.n41 avss.t248 10.5285
R2268 avss.n42 avss.t60 10.5285
R2269 avss.n43 avss.t204 10.5285
R2270 avss.n44 avss.t137 10.5285
R2271 avss.n45 avss.t210 10.5285
R2272 avss.n46 avss.t11 10.5285
R2273 avss.n47 avss.t38 10.5285
R2274 avss.n48 avss.t253 10.5285
R2275 avss.n49 avss.t28 10.5285
R2276 avss.n50 avss.t48 10.5285
R2277 avss.n51 avss.t121 10.5285
R2278 avss.n52 avss.t133 10.5285
R2279 avss.n54 avss.t65 10.5285
R2280 avss.n56 avss.t217 10.5285
R2281 avss.n104 avss.t17 10.5285
R2282 avss.n103 avss.t174 10.5285
R2283 avss.n102 avss.t83 10.5285
R2284 avss.n101 avss.t257 10.5285
R2285 avss.n100 avss.t89 10.5285
R2286 avss.n99 avss.t103 10.5285
R2287 avss.n98 avss.t234 10.5285
R2288 avss.n97 avss.t194 10.5285
R2289 avss.n96 avss.t54 10.5285
R2290 avss.n95 avss.t21 10.5285
R2291 avss.n94 avss.t96 10.5285
R2292 avss.n93 avss.t26 10.5285
R2293 avss.n92 avss.t202 10.5285
R2294 avss.n91 avss.t163 10.5285
R2295 avss.n90 avss.t141 10.5285
R2296 avss.n89 avss.t179 10.5285
R2297 avss.n88 avss.t232 10.5285
R2298 avss.n87 avss.t243 10.5285
R2299 avss.n86 avss.t42 10.5285
R2300 avss.n85 avss.t190 10.5285
R2301 avss.n84 avss.t32 10.5285
R2302 avss.n83 avss.t46 10.5285
R2303 avss.n82 avss.t154 10.5285
R2304 avss.n81 avss.t192 10.5285
R2305 avss.n80 avss.t245 10.5285
R2306 avss.n79 avss.t117 10.5285
R2307 avss.n78 avss.t113 10.5285
R2308 avss.n77 avss.t225 10.5285
R2309 avss.n76 avss.t81 10.5285
R2310 avss.n75 avss.t67 10.5285
R2311 avss.n74 avss.t159 10.5285
R2312 avss.n73 avss.t85 10.5285
R2313 avss.n72 avss.t148 10.5285
R2314 avss.n71 avss.t34 10.5285
R2315 avss.n70 avss.t220 10.5285
R2316 avss.n69 avss.t57 10.5285
R2317 avss.n68 avss.t77 10.5285
R2318 avss.n67 avss.t9 10.5285
R2319 avss.n66 avss.t151 10.5285
R2320 avss.n65 avss.t172 10.5285
R2321 avss.n64 avss.t50 10.5285
R2322 avss.n63 avss.t30 10.5285
R2323 avss.n62 avss.t251 10.5285
R2324 avss.n61 avss.t52 10.5285
R2325 avss.n60 avss.t241 10.5285
R2326 avss.n59 avss.t44 10.5285
R2327 avss.n58 avss.t198 10.5285
R2328 avss.n2 avss.t87 10.5285
R2329 avss.n0 avss.t75 10.5285
R2330 avss.n108 avss.t238 10.5285
R2331 avss.n106 avss.t109 10.5285
R2332 avss.n592 avss.n591 10.3069
R2333 avss.n605 avss.n604 7.9365
R2334 avss.n727 avss.n726 7.29749
R2335 avss.n606 avss.n258 7.2709
R2336 avss.n604 avss.n261 6.4005
R2337 avss.n588 avss.n116 5.91288
R2338 avss.n727 avss.n111 5.86875
R2339 avss.n720 avss.n127 5.34317
R2340 avss.n598 avss.n258 5.1205
R2341 avss.n721 avss.n126 3.60826
R2342 avss.n723 avss.n124 3.46074
R2343 avss.n722 avss.n125 3.42275
R2344 avss.n736 avss.n735 2.91095
R2345 avss.n735 avss.t2 2.91095
R2346 avss.n734 avss.n733 2.91095
R2347 avss.t2 avss.n734 2.91095
R2348 avss.n652 avss 2.78541
R2349 avss.n208 avss 2.23541
R2350 avss.n641 avss 2.23541
R2351 avss.n720 avss.n719 2.20222
R2352 avss.n732 avss.n113 2.19151
R2353 avss.n120 avss.n113 2.19151
R2354 avss.n114 avss.n112 2.19151
R2355 avss.t98 avss.n272 1.84498
R2356 avss.n726 avss.n122 1.80664
R2357 avss.n607 avss.n606 1.5505
R2358 avss.n609 avss.n608 1.5505
R2359 avss.n413 avss.n412 1.5505
R2360 avss.n415 avss.n414 1.5505
R2361 avss.n403 avss.n402 1.5505
R2362 avss.n393 avss.n392 1.5505
R2363 avss.n577 avss.n576 1.5505
R2364 avss.n579 avss.n578 1.5505
R2365 avss.n305 avss.n304 1.5505
R2366 avss.n618 avss.n617 1.5505
R2367 avss.n620 avss.n619 1.5505
R2368 avss.n424 avss.n423 1.5505
R2369 avss.n426 avss.n425 1.5505
R2370 avss.n564 avss.n563 1.5505
R2371 avss.n566 avss.n565 1.5505
R2372 avss.n455 avss.n454 1.5505
R2373 avss.n481 avss.n480 1.5505
R2374 avss.n550 avss.n549 1.5505
R2375 avss.n552 avss.n551 1.5505
R2376 avss.n508 avss.n507 1.5505
R2377 avss.n495 avss.n494 1.5505
R2378 avss.n284 avss.n126 1.5505
R2379 avss.n631 avss.n630 1.5505
R2380 avss.n629 avss.n628 1.5505
R2381 avss.n519 avss.n518 1.5505
R2382 avss.n197 avss.n185 1.5505
R2383 avss.n209 avss.n208 1.5505
R2384 avss.n220 avss.n127 1.5505
R2385 avss.n641 avss.n640 1.5505
R2386 avss.n53 avss.n52 1.42736
R2387 avss.n55 avss.n54 1.42736
R2388 avss.n57 avss.n56 1.42736
R2389 avss.n2 avss.n1 1.42736
R2390 avss.n108 avss.n107 1.42736
R2391 avss.n706 avss.n705 1.37676
R2392 avss.n110 avss 1.34985
R2393 avss.n705 avss.n128 1.25238
R2394 avss.n719 avss.n128 1.25238
R2395 avss avss.n577 1.23541
R2396 avss.n393 avss 1.23541
R2397 avss.n403 avss 1.23541
R2398 avss.n414 avss 1.23541
R2399 avss avss.n413 1.23541
R2400 avss.n608 avss 1.23541
R2401 avss.n565 avss 1.23541
R2402 avss avss.n564 1.23541
R2403 avss.n425 avss 1.23541
R2404 avss avss.n424 1.23541
R2405 avss.n619 avss 1.23541
R2406 avss avss.n618 1.23541
R2407 avss.n480 avss 1.23541
R2408 avss.n495 avss 1.23541
R2409 avss.n508 avss 1.23541
R2410 avss.n551 avss 1.23541
R2411 avss avss.n550 1.23541
R2412 avss.n629 avss 1.23541
R2413 avss.n630 avss 1.23541
R2414 avss avss.n126 1.23541
R2415 avss.n208 avss 1.23541
R2416 avss avss.n185 1.23541
R2417 avss avss.n127 1.23541
R2418 avss.n605 avss.n124 1.163
R2419 avss.n351 avss.n350 1.163
R2420 avss.n298 avss.n125 1.163
R2421 avss.n469 avss.n456 1.163
R2422 avss.n540 avss.n520 1.163
R2423 avss.n643 avss.n642 1.163
R2424 avss avss.n519 1.11353
R2425 avss avss.n641 1.11353
R2426 avss avss.n607 1.10745
R2427 avss.n304 avss 1.07104
R2428 avss.n726 avss.n725 0.816777
R2429 avss.n578 avss.n351 0.74738
R2430 avss.n739 avss.n109 0.714152
R2431 avss.n739 avss.n0 0.713709
R2432 avss.n456 avss.n455 0.709387
R2433 avss.n606 avss.n605 0.6661
R2434 avss.n578 avss 0.5005
R2435 avss.n577 avss 0.5005
R2436 avss avss.n393 0.5005
R2437 avss avss.n403 0.5005
R2438 avss.n414 avss 0.5005
R2439 avss.n413 avss 0.5005
R2440 avss.n608 avss 0.5005
R2441 avss.n455 avss 0.5005
R2442 avss.n565 avss 0.5005
R2443 avss.n564 avss 0.5005
R2444 avss.n425 avss 0.5005
R2445 avss.n424 avss 0.5005
R2446 avss.n619 avss 0.5005
R2447 avss.n618 avss 0.5005
R2448 avss.n480 avss 0.5005
R2449 avss avss.n495 0.5005
R2450 avss avss.n508 0.5005
R2451 avss.n551 avss 0.5005
R2452 avss.n519 avss 0.5005
R2453 avss avss.n629 0.5005
R2454 avss.n630 avss 0.5005
R2455 avss.n740 avss.n739 0.459809
R2456 avss.n708 avss.n707 0.388
R2457 avss.n703 avss.n702 0.388
R2458 avss.n679 avss.n678 0.388
R2459 avss.n717 avss.n716 0.388
R2460 avss.n738 avss.n110 0.377227
R2461 avss.n706 avss.n146 0.329037
R2462 avss.n704 avss.n147 0.329037
R2463 avss.n677 avss.n676 0.329037
R2464 avss.n718 avss.n129 0.329037
R2465 avss.n707 avss 0.301379
R2466 avss.n703 avss 0.301379
R2467 avss.n678 avss 0.301379
R2468 avss.n717 avss 0.301379
R2469 avss.n550 avss.n520 0.274922
R2470 avss.n642 avss.n185 0.274922
R2471 avss.n707 avss.n706 0.258038
R2472 avss.n704 avss.n703 0.258038
R2473 avss.n678 avss.n677 0.258038
R2474 avss.n718 avss.n717 0.258038
R2475 avss.n54 avss.n53 0.238532
R2476 avss.n56 avss.n55 0.238532
R2477 avss.n3 avss.n2 0.238532
R2478 avss.n1 avss.n0 0.238532
R2479 avss.n109 avss.n108 0.238532
R2480 avss.n107 avss.n106 0.238532
R2481 avss.n351 avss 0.221517
R2482 avss.n724 avss.n110 0.191699
R2483 avss.n456 avss 0.183525
R2484 avss.n722 avss.n721 0.161722
R2485 avss.n721 avss.n720 0.160761
R2486 avss.n723 avss.n722 0.157495
R2487 avss.n4 avss.n3 0.151652
R2488 avss.n106 avss.n105 0.151209
R2489 avss.n52 avss.n51 0.142787
R2490 avss.n58 avss.n57 0.142344
R2491 avss.n740 avss 0.136236
R2492 avss.n724 avss.n723 0.133859
R2493 avss.n705 avss.n704 0.124872
R2494 avss.n677 avss.n128 0.124872
R2495 avss.n719 avss.n718 0.124872
R2496 avss avss.n740 0.0871641
R2497 avss.n739 avss.n738 0.0830826
R2498 avss.n708 avss.n145 0.0554356
R2499 avss.n702 avss.n148 0.0554356
R2500 avss.n679 avss.n675 0.0554356
R2501 avss.n716 avss.n130 0.0554356
R2502 avss.n51 avss.n50 0.0429147
R2503 avss.n50 avss.n49 0.0429147
R2504 avss.n49 avss.n48 0.0429147
R2505 avss.n48 avss.n47 0.0429147
R2506 avss.n47 avss.n46 0.0429147
R2507 avss.n46 avss.n45 0.0429147
R2508 avss.n45 avss.n44 0.0429147
R2509 avss.n44 avss.n43 0.0429147
R2510 avss.n43 avss.n42 0.0429147
R2511 avss.n42 avss.n41 0.0429147
R2512 avss.n41 avss.n40 0.0429147
R2513 avss.n40 avss.n39 0.0429147
R2514 avss.n39 avss.n38 0.0429147
R2515 avss.n38 avss.n37 0.0429147
R2516 avss.n37 avss.n36 0.0429147
R2517 avss.n36 avss.n35 0.0429147
R2518 avss.n35 avss.n34 0.0429147
R2519 avss.n34 avss.n33 0.0429147
R2520 avss.n33 avss.n32 0.0429147
R2521 avss.n32 avss.n31 0.0429147
R2522 avss.n31 avss.n30 0.0429147
R2523 avss.n30 avss.n29 0.0429147
R2524 avss.n29 avss.n28 0.0429147
R2525 avss.n28 avss.n27 0.0429147
R2526 avss.n27 avss.n26 0.0429147
R2527 avss.n26 avss.n25 0.0429147
R2528 avss.n25 avss.n24 0.0429147
R2529 avss.n24 avss.n23 0.0429147
R2530 avss.n23 avss.n22 0.0429147
R2531 avss.n22 avss.n21 0.0429147
R2532 avss.n21 avss.n20 0.0429147
R2533 avss.n20 avss.n19 0.0429147
R2534 avss.n19 avss.n18 0.0429147
R2535 avss.n18 avss.n17 0.0429147
R2536 avss.n17 avss.n16 0.0429147
R2537 avss.n16 avss.n15 0.0429147
R2538 avss.n15 avss.n14 0.0429147
R2539 avss.n14 avss.n13 0.0429147
R2540 avss.n13 avss.n12 0.0429147
R2541 avss.n12 avss.n11 0.0429147
R2542 avss.n11 avss.n10 0.0429147
R2543 avss.n10 avss.n9 0.0429147
R2544 avss.n9 avss.n8 0.0429147
R2545 avss.n8 avss.n7 0.0429147
R2546 avss.n7 avss.n6 0.0429147
R2547 avss.n6 avss.n5 0.0429147
R2548 avss.n59 avss.n58 0.0429147
R2549 avss.n60 avss.n59 0.0429147
R2550 avss.n61 avss.n60 0.0429147
R2551 avss.n62 avss.n61 0.0429147
R2552 avss.n63 avss.n62 0.0429147
R2553 avss.n64 avss.n63 0.0429147
R2554 avss.n65 avss.n64 0.0429147
R2555 avss.n66 avss.n65 0.0429147
R2556 avss.n67 avss.n66 0.0429147
R2557 avss.n68 avss.n67 0.0429147
R2558 avss.n69 avss.n68 0.0429147
R2559 avss.n70 avss.n69 0.0429147
R2560 avss.n71 avss.n70 0.0429147
R2561 avss.n72 avss.n71 0.0429147
R2562 avss.n73 avss.n72 0.0429147
R2563 avss.n74 avss.n73 0.0429147
R2564 avss.n75 avss.n74 0.0429147
R2565 avss.n76 avss.n75 0.0429147
R2566 avss.n77 avss.n76 0.0429147
R2567 avss.n78 avss.n77 0.0429147
R2568 avss.n79 avss.n78 0.0429147
R2569 avss.n80 avss.n79 0.0429147
R2570 avss.n81 avss.n80 0.0429147
R2571 avss.n82 avss.n81 0.0429147
R2572 avss.n83 avss.n82 0.0429147
R2573 avss.n84 avss.n83 0.0429147
R2574 avss.n85 avss.n84 0.0429147
R2575 avss.n86 avss.n85 0.0429147
R2576 avss.n87 avss.n86 0.0429147
R2577 avss.n88 avss.n87 0.0429147
R2578 avss.n89 avss.n88 0.0429147
R2579 avss.n90 avss.n89 0.0429147
R2580 avss.n91 avss.n90 0.0429147
R2581 avss.n92 avss.n91 0.0429147
R2582 avss.n93 avss.n92 0.0429147
R2583 avss.n94 avss.n93 0.0429147
R2584 avss.n95 avss.n94 0.0429147
R2585 avss.n96 avss.n95 0.0429147
R2586 avss.n97 avss.n96 0.0429147
R2587 avss.n98 avss.n97 0.0429147
R2588 avss.n99 avss.n98 0.0429147
R2589 avss.n100 avss.n99 0.0429147
R2590 avss.n101 avss.n100 0.0429147
R2591 avss.n102 avss.n101 0.0429147
R2592 avss.n103 avss.n102 0.0429147
R2593 avss.n104 avss.n103 0.0429147
R2594 avss.n520 avss 0.0390514
R2595 avss.n642 avss 0.0390514
R2596 avss.n5 avss.n4 0.0270934
R2597 avss.n105 avss.n104 0.0270934
R2598 avss.n725 avss.n724 0.025588
R2599 avss.n607 avss.n124 0.00896354
R2600 avss.n738 avss.n737 0.00821144
R2601 avss.n304 avss.n125 0.00738559
R2602 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t1 227.512
R2603 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t4 99.4875
R2604 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t2 99.1756
R2605 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t0 41.0738
R2606 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t6 22.2871
R2607 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n0 21.2032
R2608 multiplexer_0.vtrip_1_b.n0 multiplexer_0.vtrip_1_b.t9 16.8731
R2609 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t12 16.8731
R2610 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t5 16.8731
R2611 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t8 16.8731
R2612 multiplexer_0.vtrip_1_b.n0 multiplexer_0.vtrip_1_b.t10 16.5088
R2613 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t3 16.5088
R2614 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t7 16.5088
R2615 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.t11 16.5088
R2616 dvdd.n534 dvdd.n98 6151.76
R2617 dvdd.n528 dvdd.n98 6151.76
R2618 dvdd.n528 dvdd.n57 6151.76
R2619 dvdd.n546 dvdd.n57 6151.76
R2620 dvdd.n546 dvdd.n71 6151.76
R2621 dvdd.n633 dvdd.n71 6151.76
R2622 dvdd.n533 dvdd.n99 6151.76
R2623 dvdd.n527 dvdd.n99 6151.76
R2624 dvdd.n527 dvdd.n58 6151.76
R2625 dvdd.n545 dvdd.n58 6151.76
R2626 dvdd.n545 dvdd.n72 6151.76
R2627 dvdd.n635 dvdd.n72 6151.76
R2628 dvdd.n622 dvdd.n94 6151.76
R2629 dvdd.n622 dvdd.n96 6151.76
R2630 dvdd.n96 dvdd.n59 6151.76
R2631 dvdd.n543 dvdd.n59 6151.76
R2632 dvdd.n543 dvdd.n73 6151.76
R2633 dvdd.n632 dvdd.n73 6151.76
R2634 dvdd.n621 dvdd.n101 6151.76
R2635 dvdd.n621 dvdd.n53 6151.76
R2636 dvdd.n659 dvdd.n53 6151.76
R2637 dvdd.n659 dvdd.n54 6151.76
R2638 dvdd.n653 dvdd.n54 6151.76
R2639 dvdd.n653 dvdd.n74 6151.76
R2640 dvdd.n111 dvdd.n100 6151.76
R2641 dvdd.n100 dvdd.n60 6151.76
R2642 dvdd.n658 dvdd.n60 6151.76
R2643 dvdd.n658 dvdd.n61 6151.76
R2644 dvdd.n654 dvdd.n61 6151.76
R2645 dvdd.n654 dvdd.n69 6151.76
R2646 dvdd.n589 dvdd.n268 4207.06
R2647 dvdd.n592 dvdd.n591 4207.06
R2648 dvdd.n227 dvdd.n139 3328.24
R2649 dvdd.n147 dvdd.n139 3328.24
R2650 dvdd.n242 dvdd.n132 3328.24
R2651 dvdd.n243 dvdd.n242 3328.24
R2652 dvdd.n169 dvdd.n138 3328.24
R2653 dvdd.n182 dvdd.n138 3328.24
R2654 dvdd.n201 dvdd.n137 3328.24
R2655 dvdd.n191 dvdd.n137 3328.24
R2656 dvdd.n170 dvdd.n136 3328.24
R2657 dvdd.n193 dvdd.n136 3328.24
R2658 dvdd.n241 dvdd.n141 3328.24
R2659 dvdd.n241 dvdd.n142 3328.24
R2660 dvdd.n216 dvdd.n140 3328.24
R2661 dvdd.n236 dvdd.n140 3328.24
R2662 dvdd.n562 dvdd.n557 2822.48
R2663 dvdd.n560 dvdd.n559 2822.48
R2664 dvdd.n596 dvdd.n263 2442.35
R2665 dvdd.n599 dvdd.n262 2442.35
R2666 dvdd.n569 dvdd.n554 2442.35
R2667 dvdd.n576 dvdd.n519 2442.35
R2668 dvdd.n584 dvdd.n583 2442.35
R2669 dvdd.n581 dvdd.n274 2442.35
R2670 dvdd.n44 dvdd.n43 2442.35
R2671 dvdd.n41 dvdd.n39 2442.35
R2672 dvdd.n32 dvdd.n31 2442.35
R2673 dvdd.n29 dvdd.n27 2442.35
R2674 dvdd.n20 dvdd.n19 2442.35
R2675 dvdd.n17 dvdd.n15 2442.35
R2676 dvdd.n8 dvdd.n7 2442.35
R2677 dvdd.n5 dvdd.n3 2442.35
R2678 dvdd.n194 dvdd.n122 1736.47
R2679 dvdd.n175 dvdd.n155 1736.47
R2680 dvdd.n225 dvdd.n160 1736.47
R2681 dvdd.n254 dvdd.n124 1736.47
R2682 dvdd.n602 dvdd.n106 1736.47
R2683 dvdd.n86 dvdd.n80 1736.47
R2684 dvdd.n617 dvdd.n104 1736.47
R2685 dvdd.n649 dvdd.n78 1736.47
R2686 dvdd.n574 dvdd.n522 1563.53
R2687 dvdd.n569 dvdd.n522 1563.53
R2688 dvdd.n576 dvdd.n520 1563.53
R2689 dvdd.n567 dvdd.n520 1563.53
R2690 dvdd.n268 dvdd.n266 1068.61
R2691 dvdd.n591 dvdd.n590 1068.61
R2692 dvdd.n201 dvdd.n200 878.823
R2693 dvdd.n200 dvdd.n170 878.823
R2694 dvdd.n173 dvdd.n163 878.823
R2695 dvdd.n174 dvdd.n173 878.823
R2696 dvdd.n202 dvdd.n169 878.823
R2697 dvdd.n202 dvdd.n201 878.823
R2698 dvdd.n145 dvdd.n123 878.823
R2699 dvdd.n244 dvdd.n123 878.823
R2700 dvdd.n209 dvdd.n208 878.823
R2701 dvdd.n208 dvdd.n163 878.823
R2702 dvdd.n168 dvdd.n132 878.823
R2703 dvdd.n169 dvdd.n168 878.823
R2704 dvdd.n236 dvdd.n234 878.823
R2705 dvdd.n234 dvdd.n147 878.823
R2706 dvdd.n214 dvdd.n213 878.823
R2707 dvdd.n214 dvdd.n153 878.823
R2708 dvdd.n210 dvdd.n153 878.823
R2709 dvdd.n210 dvdd.n209 878.823
R2710 dvdd.n216 dvdd.n152 878.823
R2711 dvdd.n227 dvdd.n152 878.823
R2712 dvdd.n228 dvdd.n227 878.823
R2713 dvdd.n228 dvdd.n132 878.823
R2714 dvdd.n147 dvdd.n130 878.823
R2715 dvdd.n243 dvdd.n130 878.823
R2716 dvdd.n243 dvdd.n131 878.823
R2717 dvdd.n182 dvdd.n131 878.823
R2718 dvdd.n244 dvdd.n121 878.823
R2719 dvdd.n121 dvdd.n118 878.823
R2720 dvdd.n256 dvdd.n118 878.823
R2721 dvdd.n256 dvdd.n119 878.823
R2722 dvdd.n182 dvdd.n180 878.823
R2723 dvdd.n191 dvdd.n180 878.823
R2724 dvdd.n192 dvdd.n191 878.823
R2725 dvdd.n193 dvdd.n192 878.823
R2726 dvdd.n122 dvdd.n119 878.823
R2727 dvdd.n175 dvdd.n174 878.823
R2728 dvdd.n237 dvdd.n142 878.823
R2729 dvdd.n237 dvdd.n236 878.823
R2730 dvdd.n217 dvdd.n141 878.823
R2731 dvdd.n217 dvdd.n216 878.823
R2732 dvdd.n254 dvdd.n125 878.823
R2733 dvdd.n125 dvdd.n120 878.823
R2734 dvdd.n145 dvdd.n120 878.823
R2735 dvdd.n213 dvdd.n160 878.823
R2736 dvdd.n65 dvdd.n54 878.823
R2737 dvdd.n65 dvdd.n61 878.823
R2738 dvdd.n608 dvdd.n109 878.823
R2739 dvdd.n608 dvdd.n607 878.823
R2740 dvdd.n611 dvdd.n111 878.823
R2741 dvdd.n611 dvdd.n94 878.823
R2742 dvdd.n95 dvdd.n60 878.823
R2743 dvdd.n96 dvdd.n95 878.823
R2744 dvdd.n542 dvdd.n61 878.823
R2745 dvdd.n543 dvdd.n542 878.823
R2746 dvdd.n607 dvdd.n606 878.823
R2747 dvdd.n606 dvdd.n115 878.823
R2748 dvdd.n532 dvdd.n94 878.823
R2749 dvdd.n533 dvdd.n532 878.823
R2750 dvdd.n526 dvdd.n96 878.823
R2751 dvdd.n527 dvdd.n526 878.823
R2752 dvdd.n544 dvdd.n543 878.823
R2753 dvdd.n545 dvdd.n544 878.823
R2754 dvdd.n602 dvdd.n115 878.823
R2755 dvdd.n535 dvdd.n533 878.823
R2756 dvdd.n535 dvdd.n534 878.823
R2757 dvdd.n529 dvdd.n527 878.823
R2758 dvdd.n529 dvdd.n528 878.823
R2759 dvdd.n547 dvdd.n545 878.823
R2760 dvdd.n547 dvdd.n546 878.823
R2761 dvdd.n86 dvdd.n85 878.823
R2762 dvdd.n636 dvdd.n632 878.823
R2763 dvdd.n636 dvdd.n635 878.823
R2764 dvdd.n635 dvdd.n634 878.823
R2765 dvdd.n634 dvdd.n633 878.823
R2766 dvdd.n644 dvdd.n83 878.823
R2767 dvdd.n644 dvdd.n643 878.823
R2768 dvdd.n643 dvdd.n642 878.823
R2769 dvdd.n642 dvdd.n85 878.823
R2770 dvdd.n62 dvdd.n53 878.823
R2771 dvdd.n62 dvdd.n60 878.823
R2772 dvdd.n110 dvdd.n101 878.823
R2773 dvdd.n111 dvdd.n110 878.823
R2774 dvdd.n109 dvdd.n104 878.823
R2775 dvdd.n75 dvdd.n74 878.823
R2776 dvdd.n75 dvdd.n69 878.823
R2777 dvdd.n631 dvdd.n69 878.823
R2778 dvdd.n632 dvdd.n631 878.823
R2779 dvdd.n83 dvdd.n78 878.823
R2780 dvdd.n524 dvdd.n522 878.823
R2781 dvdd.n524 dvdd.n520 878.823
R2782 dvdd.n226 dvdd.n153 857.648
R2783 dvdd.n227 dvdd.n226 857.648
R2784 dvdd.n147 dvdd.n146 857.648
R2785 dvdd.n146 dvdd.n145 857.648
R2786 dvdd.n209 dvdd.n158 857.648
R2787 dvdd.n158 dvdd.n132 857.648
R2788 dvdd.n245 dvdd.n243 857.648
R2789 dvdd.n245 dvdd.n244 857.648
R2790 dvdd.n163 dvdd.n157 857.648
R2791 dvdd.n169 dvdd.n157 857.648
R2792 dvdd.n183 dvdd.n182 857.648
R2793 dvdd.n183 dvdd.n118 857.648
R2794 dvdd.n174 dvdd.n156 857.648
R2795 dvdd.n201 dvdd.n156 857.648
R2796 dvdd.n191 dvdd.n190 857.648
R2797 dvdd.n190 dvdd.n119 857.648
R2798 dvdd.n170 dvdd.n155 857.648
R2799 dvdd.n194 dvdd.n193 857.648
R2800 dvdd.n225 dvdd.n141 857.648
R2801 dvdd.n142 dvdd.n124 857.648
R2802 dvdd.n213 dvdd.n159 857.648
R2803 dvdd.n216 dvdd.n159 857.648
R2804 dvdd.n236 dvdd.n235 857.648
R2805 dvdd.n235 dvdd.n125 857.648
R2806 dvdd.n534 dvdd.n106 857.648
R2807 dvdd.n633 dvdd.n80 857.648
R2808 dvdd.n115 dvdd.n107 857.648
R2809 dvdd.n533 dvdd.n107 857.648
R2810 dvdd.n635 dvdd.n81 857.648
R2811 dvdd.n85 dvdd.n81 857.648
R2812 dvdd.n607 dvdd.n108 857.648
R2813 dvdd.n108 dvdd.n94 857.648
R2814 dvdd.n632 dvdd.n82 857.648
R2815 dvdd.n643 dvdd.n82 857.648
R2816 dvdd.n617 dvdd.n101 857.648
R2817 dvdd.n649 dvdd.n74 857.648
R2818 dvdd.n616 dvdd.n109 857.648
R2819 dvdd.n616 dvdd.n111 857.648
R2820 dvdd.n648 dvdd.n69 857.648
R2821 dvdd.n648 dvdd.n83 857.648
R2822 dvdd.t15 dvdd.n97 741.205
R2823 dvdd.t15 dvdd.n55 741.205
R2824 dvdd.t26 dvdd.n55 741.205
R2825 dvdd.t26 dvdd.n56 741.205
R2826 dvdd.t44 dvdd.n56 741.205
R2827 dvdd.t44 dvdd.n70 741.205
R2828 dvdd.t119 dvdd.n521 659.64
R2829 dvdd.t94 dvdd.n521 659.64
R2830 dvdd.n552 dvdd.n551 656.188
R2831 dvdd.n551 dvdd.n550 656.188
R2832 dvdd.n538 dvdd.n537 656.188
R2833 dvdd.n539 dvdd.n538 656.188
R2834 dvdd.n540 dvdd.n539 656.188
R2835 dvdd.n541 dvdd.n540 656.188
R2836 dvdd.n541 dvdd.n89 656.188
R2837 dvdd.n638 dvdd.n89 656.188
R2838 dvdd.n623 dvdd.n93 656.188
R2839 dvdd.n624 dvdd.n623 656.188
R2840 dvdd.n625 dvdd.n624 656.188
R2841 dvdd.n626 dvdd.n625 656.188
R2842 dvdd.n627 dvdd.n626 656.188
R2843 dvdd.n629 dvdd.n627 656.188
R2844 dvdd.n614 dvdd.n613 656.188
R2845 dvdd.n613 dvdd.n64 656.188
R2846 dvdd.n657 dvdd.n64 656.188
R2847 dvdd.n657 dvdd.n656 656.188
R2848 dvdd.n656 dvdd.n655 656.188
R2849 dvdd.n655 dvdd.n68 656.188
R2850 dvdd.n563 dvdd.n556 545.13
R2851 dvdd.n556 dvdd.n275 545.13
R2852 dvdd.n575 dvdd.n519 535.419
R2853 dvdd.n568 dvdd.n554 535.419
R2854 dvdd.n274 dvdd.n272 535.419
R2855 dvdd.n583 dvdd.n582 535.419
R2856 dvdd.n39 dvdd.n38 535.419
R2857 dvdd.n43 dvdd.n42 535.419
R2858 dvdd.n27 dvdd.n26 535.419
R2859 dvdd.n31 dvdd.n30 535.419
R2860 dvdd.n15 dvdd.n14 535.419
R2861 dvdd.n19 dvdd.n18 535.419
R2862 dvdd.n3 dvdd.n2 535.419
R2863 dvdd.n7 dvdd.n6 535.419
R2864 dvdd.n553 dvdd.n552 436.104
R2865 dvdd.n240 dvdd.n143 355.012
R2866 dvdd.n240 dvdd.n239 355.012
R2867 dvdd.n220 dvdd.n219 355.012
R2868 dvdd.n219 dvdd.n144 355.012
R2869 dvdd.n231 dvdd.n230 355.012
R2870 dvdd.n232 dvdd.n231 355.012
R2871 dvdd.n151 dvdd.n133 355.012
R2872 dvdd.n133 dvdd.n129 355.012
R2873 dvdd.n204 dvdd.n166 355.012
R2874 dvdd.n185 dvdd.n166 355.012
R2875 dvdd.n187 dvdd.n167 355.012
R2876 dvdd.n188 dvdd.n187 355.012
R2877 dvdd.n198 dvdd.n197 355.012
R2878 dvdd.n197 dvdd.n196 355.012
R2879 dvdd.n594 dvdd.n593 348.613
R2880 dvdd.n593 dvdd.n265 348.613
R2881 dvdd.n559 dvdd.n558 318.108
R2882 dvdd.n562 dvdd.n561 318.108
R2883 dvdd.n565 dvdd.n563 295.529
R2884 dvdd.n578 dvdd.n275 295.529
R2885 dvdd.t1 dvdd.n134 271.635
R2886 dvdd.t1 dvdd.n135 271.635
R2887 dvdd.n40 dvdd.n36 260.519
R2888 dvdd.n28 dvdd.n24 260.519
R2889 dvdd.n16 dvdd.n12 260.519
R2890 dvdd.n4 dvdd.n0 260.519
R2891 dvdd.n600 dvdd.n261 260.329
R2892 dvdd.n601 dvdd.n600 243.018
R2893 dvdd.n594 dvdd.n261 229.702
R2894 dvdd.n422 dvdd.t98 229.419
R2895 dvdd.n477 dvdd.t102 229.419
R2896 dvdd.n48 dvdd.t101 229.419
R2897 dvdd.n508 dvdd.t120 229.212
R2898 dvdd.n505 dvdd.t117 229.212
R2899 dvdd.n507 dvdd.t107 229.179
R2900 dvdd.n417 dvdd.t118 229.076
R2901 dvdd.n47 dvdd.t93 228.484
R2902 dvdd.n35 dvdd.t112 228.484
R2903 dvdd.n23 dvdd.t110 228.484
R2904 dvdd.n11 dvdd.t97 228.484
R2905 dvdd.n422 dvdd.t103 228.215
R2906 dvdd.n298 dvdd.t52 228.215
R2907 dvdd.n419 dvdd.t113 228.215
R2908 dvdd.n418 dvdd.t114 228.215
R2909 dvdd.n417 dvdd.t115 228.215
R2910 dvdd.n294 dvdd.t61 228.215
R2911 dvdd.n495 dvdd.t76 228.215
R2912 dvdd.n398 dvdd.t31 228.215
R2913 dvdd.n283 dvdd.t16 228.215
R2914 dvdd.n510 dvdd.t27 228.215
R2915 dvdd.n514 dvdd.t28 228.215
R2916 dvdd.n517 dvdd.t95 228.215
R2917 dvdd.n278 dvdd.t45 228.215
R2918 dvdd.n452 dvdd.t24 228.215
R2919 dvdd.n454 dvdd.t23 228.215
R2920 dvdd.n450 dvdd.t20 228.215
R2921 dvdd.n448 dvdd.t21 228.215
R2922 dvdd.n446 dvdd.t72 228.215
R2923 dvdd.n444 dvdd.t73 228.215
R2924 dvdd.n435 dvdd.t54 228.215
R2925 dvdd.n433 dvdd.t55 228.215
R2926 dvdd.n477 dvdd.t105 228.215
R2927 dvdd.n48 dvdd.t104 228.215
R2928 dvdd.n431 dvdd.t58 228.215
R2929 dvdd.n428 dvdd.t57 228.215
R2930 dvdd.n436 dvdd.t67 228.215
R2931 dvdd.n437 dvdd.t66 228.215
R2932 dvdd.n455 dvdd.t46 228.215
R2933 dvdd.n281 dvdd.t17 228.215
R2934 dvdd.n383 dvdd.t85 228.215
R2935 dvdd.n319 dvdd.t84 228.215
R2936 dvdd.n318 dvdd.t81 228.215
R2937 dvdd.n313 dvdd.t12 228.215
R2938 dvdd.n311 dvdd.t13 228.215
R2939 dvdd.n309 dvdd.t9 228.215
R2940 dvdd.n307 dvdd.t10 228.215
R2941 dvdd.n305 dvdd.t6 228.215
R2942 dvdd.n303 dvdd.t7 228.215
R2943 dvdd.n301 dvdd.t78 228.215
R2944 dvdd.n351 dvdd.t38 228.215
R2945 dvdd.n344 dvdd.t63 228.215
R2946 dvdd.n340 dvdd.t69 228.215
R2947 dvdd.n336 dvdd.t87 228.215
R2948 dvdd.n332 dvdd.t41 228.215
R2949 dvdd.n323 dvdd.t2 228.215
R2950 dvdd.n321 dvdd.t3 228.215
R2951 dvdd.n329 dvdd.t48 228.215
R2952 dvdd.n324 dvdd.t49 228.215
R2953 dvdd.n326 dvdd.t42 228.215
R2954 dvdd.n334 dvdd.t88 228.215
R2955 dvdd.n338 dvdd.t70 228.215
R2956 dvdd.n342 dvdd.t64 228.215
R2957 dvdd.n346 dvdd.t39 228.215
R2958 dvdd.n348 dvdd.t90 228.215
R2959 dvdd.n355 dvdd.t91 228.215
R2960 dvdd.n299 dvdd.t79 228.215
R2961 dvdd.n397 dvdd.t82 228.215
R2962 dvdd.n385 dvdd.t34 228.215
R2963 dvdd.n284 dvdd.t35 228.215
R2964 dvdd.n286 dvdd.t32 228.215
R2965 dvdd.n291 dvdd.t75 228.215
R2966 dvdd.n292 dvdd.t60 228.215
R2967 dvdd.n295 dvdd.t51 228.215
R2968 dvdd.n597 dvdd.n596 214.912
R2969 dvdd.n599 dvdd.n598 214.912
R2970 dvdd.n177 dvdd.n176 185.225
R2971 dvdd.n224 dvdd.n223 185.225
R2972 dvdd.n549 dvdd.n87 185.225
R2973 dvdd.n40 dvdd.n37 176.139
R2974 dvdd.n28 dvdd.n25 176.139
R2975 dvdd.n16 dvdd.n13 176.139
R2976 dvdd.n4 dvdd.n1 176.139
R2977 dvdd.n603 dvdd.n601 167.906
R2978 dvdd.n580 dvdd.n265 160.376
R2979 dvdd.n580 dvdd.n579 160.376
R2980 dvdd.t59 dvdd.n489 120.174
R2981 dvdd.n490 dvdd.t59 120.174
R2982 dvdd.n493 dvdd.t74 120.174
R2983 dvdd.t74 dvdd.n289 120.174
R2984 dvdd.n462 dvdd.t22 120.174
R2985 dvdd.t22 dvdd.n461 120.174
R2986 dvdd.t18 dvdd.n465 120.174
R2987 dvdd.n466 dvdd.t18 120.174
R2988 dvdd.t71 dvdd.n469 120.174
R2989 dvdd.n470 dvdd.t71 120.174
R2990 dvdd.t53 dvdd.n473 120.174
R2991 dvdd.n474 dvdd.t53 120.174
R2992 dvdd.t33 dvdd.n285 120.174
R2993 dvdd.n388 dvdd.t33 120.174
R2994 dvdd.t83 dvdd.n391 120.174
R2995 dvdd.n392 dvdd.t83 120.174
R2996 dvdd.t8 dvdd.n406 120.174
R2997 dvdd.n407 dvdd.t8 120.174
R2998 dvdd.t4 dvdd.n410 120.174
R2999 dvdd.n411 dvdd.t4 120.174
R3000 dvdd.t77 dvdd.n414 120.174
R3001 dvdd.n415 dvdd.t77 120.174
R3002 dvdd.n352 dvdd.t36 120.174
R3003 dvdd.t36 dvdd.n347 120.174
R3004 dvdd.t62 dvdd.n362 120.174
R3005 dvdd.n363 dvdd.t62 120.174
R3006 dvdd.t68 dvdd.n366 120.174
R3007 dvdd.n367 dvdd.t68 120.174
R3008 dvdd.t86 dvdd.n370 120.174
R3009 dvdd.n371 dvdd.t86 120.174
R3010 dvdd.t40 dvdd.n374 120.174
R3011 dvdd.n375 dvdd.t40 120.174
R3012 dvdd.t47 dvdd.n325 120.174
R3013 dvdd.n328 dvdd.t47 120.174
R3014 dvdd.n403 dvdd.t11 120.174
R3015 dvdd.t11 dvdd.n402 120.174
R3016 dvdd.t80 dvdd.n315 120.174
R3017 dvdd.n395 dvdd.t80 120.174
R3018 dvdd.n499 dvdd.t29 120.174
R3019 dvdd.t29 dvdd.n498 120.174
R3020 dvdd.n46 dvdd.n36 118.127
R3021 dvdd.n34 dvdd.n24 118.127
R3022 dvdd.n22 dvdd.n12 118.127
R3023 dvdd.n10 dvdd.n0 118.127
R3024 dvdd.t30 dvdd.n105 103.335
R3025 dvdd.t30 dvdd.n97 103.335
R3026 dvdd.t19 dvdd.n70 103.335
R3027 dvdd.t19 dvdd.n79 103.335
R3028 dvdd.n610 dvdd.n112 100.141
R3029 dvdd.n610 dvdd.n609 100.141
R3030 dvdd.n609 dvdd.n114 100.141
R3031 dvdd.n605 dvdd.n604 100.141
R3032 dvdd.n604 dvdd.n603 100.141
R3033 dvdd.n536 dvdd.n270 98.7449
R3034 dvdd.n650 dvdd.n77 96.5745
R3035 dvdd.n222 dvdd.n215 93.7417
R3036 dvdd.n215 dvdd.n212 93.7417
R3037 dvdd.n212 dvdd.n211 93.7417
R3038 dvdd.n211 dvdd.n162 93.7417
R3039 dvdd.n207 dvdd.n162 93.7417
R3040 dvdd.n207 dvdd.n206 93.7417
R3041 dvdd.n206 dvdd.n164 93.7417
R3042 dvdd.n172 dvdd.n164 93.7417
R3043 dvdd.n176 dvdd.n172 93.7417
R3044 dvdd.n239 dvdd.n238 93.7417
R3045 dvdd.n238 dvdd.n144 93.7417
R3046 dvdd.n223 dvdd.n222 93.7417
R3047 dvdd.n218 dvdd.n143 93.7417
R3048 dvdd.n220 dvdd.n218 93.7417
R3049 dvdd.n220 dvdd.n149 93.7417
R3050 dvdd.n230 dvdd.n149 93.7417
R3051 dvdd.n233 dvdd.n144 93.7417
R3052 dvdd.n233 dvdd.n232 93.7417
R3053 dvdd.n232 dvdd.n148 93.7417
R3054 dvdd.n148 dvdd.n129 93.7417
R3055 dvdd.n230 dvdd.n229 93.7417
R3056 dvdd.n229 dvdd.n151 93.7417
R3057 dvdd.n165 dvdd.n151 93.7417
R3058 dvdd.n204 dvdd.n165 93.7417
R3059 dvdd.n181 dvdd.n129 93.7417
R3060 dvdd.n185 dvdd.n181 93.7417
R3061 dvdd.n186 dvdd.n185 93.7417
R3062 dvdd.n188 dvdd.n186 93.7417
R3063 dvdd.n204 dvdd.n203 93.7417
R3064 dvdd.n203 dvdd.n167 93.7417
R3065 dvdd.n199 dvdd.n167 93.7417
R3066 dvdd.n199 dvdd.n198 93.7417
R3067 dvdd.n188 dvdd.n178 93.7417
R3068 dvdd.n196 dvdd.n178 93.7417
R3069 dvdd.n651 dvdd.n76 93.7417
R3070 dvdd.n76 dvdd.n68 93.7417
R3071 dvdd.n66 dvdd.n52 93.7417
R3072 dvdd.n656 dvdd.n66 93.7417
R3073 dvdd.n614 dvdd.n612 93.7417
R3074 dvdd.n612 dvdd.n93 93.7417
R3075 dvdd.n91 dvdd.n64 93.7417
R3076 dvdd.n624 dvdd.n91 93.7417
R3077 dvdd.n656 dvdd.n67 93.7417
R3078 dvdd.n626 dvdd.n67 93.7417
R3079 dvdd.n531 dvdd.n93 93.7417
R3080 dvdd.n537 dvdd.n531 93.7417
R3081 dvdd.n537 dvdd.n536 93.7417
R3082 dvdd.n624 dvdd.n92 93.7417
R3083 dvdd.n539 dvdd.n92 93.7417
R3084 dvdd.n539 dvdd.n530 93.7417
R3085 dvdd.n530 dvdd.n271 93.7417
R3086 dvdd.n626 dvdd.n90 93.7417
R3087 dvdd.n541 dvdd.n90 93.7417
R3088 dvdd.n548 dvdd.n541 93.7417
R3089 dvdd.n552 dvdd.n548 93.7417
R3090 dvdd.n638 dvdd.n88 93.7417
R3091 dvdd.n550 dvdd.n88 93.7417
R3092 dvdd.n641 dvdd.n84 93.7417
R3093 dvdd.n641 dvdd.n640 93.7417
R3094 dvdd.n640 dvdd.n87 93.7417
R3095 dvdd.n630 dvdd.n68 93.7417
R3096 dvdd.n630 dvdd.n629 93.7417
R3097 dvdd.n637 dvdd.n629 93.7417
R3098 dvdd.n638 dvdd.n637 93.7417
R3099 dvdd.n63 dvdd.n51 93.7417
R3100 dvdd.n64 dvdd.n63 93.7417
R3101 dvdd.n646 dvdd.n77 93.7417
R3102 dvdd.n646 dvdd.n645 93.7417
R3103 dvdd.n645 dvdd.n84 93.7417
R3104 dvdd.n619 dvdd.n102 93.7417
R3105 dvdd.n614 dvdd.n102 93.7417
R3106 dvdd.n112 dvdd.n103 93.7417
R3107 dvdd.n605 dvdd.n258 93.7417
R3108 dvdd.n572 dvdd.n525 93.7417
R3109 dvdd.n555 dvdd.n525 93.7417
R3110 dvdd.n253 dvdd.n126 91.6685
R3111 dvdd.n195 dvdd.n179 91.6685
R3112 dvdd.n224 dvdd.n143 91.4829
R3113 dvdd.n239 dvdd.n126 91.4829
R3114 dvdd.n222 dvdd.n221 91.4829
R3115 dvdd.n221 dvdd.n220 91.4829
R3116 dvdd.n144 dvdd.n127 91.4829
R3117 dvdd.n212 dvdd.n150 91.4829
R3118 dvdd.n230 dvdd.n150 91.4829
R3119 dvdd.n232 dvdd.n128 91.4829
R3120 dvdd.n162 dvdd.n161 91.4829
R3121 dvdd.n161 dvdd.n151 91.4829
R3122 dvdd.n246 dvdd.n129 91.4829
R3123 dvdd.n206 dvdd.n205 91.4829
R3124 dvdd.n205 dvdd.n204 91.4829
R3125 dvdd.n185 dvdd.n184 91.4829
R3126 dvdd.n172 dvdd.n171 91.4829
R3127 dvdd.n171 dvdd.n167 91.4829
R3128 dvdd.n189 dvdd.n188 91.4829
R3129 dvdd.n198 dvdd.n177 91.4829
R3130 dvdd.n196 dvdd.n195 91.4829
R3131 dvdd.n550 dvdd.n549 91.4829
R3132 dvdd.n537 dvdd.n259 91.4829
R3133 dvdd.n639 dvdd.n638 91.4829
R3134 dvdd.n640 dvdd.n639 91.4829
R3135 dvdd.n113 dvdd.n93 91.4829
R3136 dvdd.n629 dvdd.n628 91.4829
R3137 dvdd.n628 dvdd.n84 91.4829
R3138 dvdd.n615 dvdd.n614 91.4829
R3139 dvdd.n647 dvdd.n68 91.4829
R3140 dvdd.n647 dvdd.n646 91.4829
R3141 dvdd.n252 dvdd.n127 85.0829
R3142 dvdd.n250 dvdd.n128 85.0829
R3143 dvdd.n248 dvdd.n246 85.0829
R3144 dvdd.n184 dvdd.n116 85.0829
R3145 dvdd.n189 dvdd.n117 85.0829
R3146 dvdd.n604 dvdd.n259 85.0829
R3147 dvdd.n114 dvdd.n113 85.0829
R3148 dvdd.n615 dvdd.n610 85.0829
R3149 dvdd.n386 dvdd.t100 84.9815
R3150 dvdd.t37 dvdd.n154 69.9975
R3151 dvdd.t37 dvdd.n134 69.9975
R3152 dvdd.n135 dvdd.t5 69.9975
R3153 dvdd.n255 dvdd.t5 69.9975
R3154 dvdd.n579 dvdd.n578 44.796
R3155 dvdd.n45 dvdd.n37 44.2181
R3156 dvdd.n33 dvdd.n25 44.2181
R3157 dvdd.n21 dvdd.n13 44.2181
R3158 dvdd.n9 dvdd.n1 44.2181
R3159 dvdd.n565 dvdd.n564 38.4243
R3160 dvdd.n225 dvdd.n224 37.0005
R3161 dvdd.t37 dvdd.n225 37.0005
R3162 dvdd.n126 dvdd.n124 37.0005
R3163 dvdd.n124 dvdd.t5 37.0005
R3164 dvdd.n221 dvdd.n159 37.0005
R3165 dvdd.t37 dvdd.n159 37.0005
R3166 dvdd.n235 dvdd.n127 37.0005
R3167 dvdd.n235 dvdd.t5 37.0005
R3168 dvdd.n226 dvdd.n150 37.0005
R3169 dvdd.n226 dvdd.t37 37.0005
R3170 dvdd.n146 dvdd.n128 37.0005
R3171 dvdd.n146 dvdd.t5 37.0005
R3172 dvdd.n161 dvdd.n158 37.0005
R3173 dvdd.t37 dvdd.n158 37.0005
R3174 dvdd.n246 dvdd.n245 37.0005
R3175 dvdd.n245 dvdd.t5 37.0005
R3176 dvdd.n205 dvdd.n157 37.0005
R3177 dvdd.t37 dvdd.n157 37.0005
R3178 dvdd.n184 dvdd.n183 37.0005
R3179 dvdd.n183 dvdd.t5 37.0005
R3180 dvdd.n171 dvdd.n156 37.0005
R3181 dvdd.t37 dvdd.n156 37.0005
R3182 dvdd.n190 dvdd.n189 37.0005
R3183 dvdd.n190 dvdd.t5 37.0005
R3184 dvdd.n195 dvdd.n194 37.0005
R3185 dvdd.n194 dvdd.t5 37.0005
R3186 dvdd.n177 dvdd.n155 37.0005
R3187 dvdd.t37 dvdd.n155 37.0005
R3188 dvdd.n262 dvdd.n260 37.0005
R3189 dvdd.n113 dvdd.n108 37.0005
R3190 dvdd.t30 dvdd.n108 37.0005
R3191 dvdd.n259 dvdd.n107 37.0005
R3192 dvdd.t30 dvdd.n107 37.0005
R3193 dvdd.n628 dvdd.n82 37.0005
R3194 dvdd.t19 dvdd.n82 37.0005
R3195 dvdd.n639 dvdd.n81 37.0005
R3196 dvdd.t19 dvdd.n81 37.0005
R3197 dvdd.n549 dvdd.n80 37.0005
R3198 dvdd.t19 dvdd.n80 37.0005
R3199 dvdd.n269 dvdd.n106 37.0005
R3200 dvdd.t30 dvdd.n106 37.0005
R3201 dvdd.n616 dvdd.n615 37.0005
R3202 dvdd.t30 dvdd.n616 37.0005
R3203 dvdd.n648 dvdd.n647 37.0005
R3204 dvdd.t19 dvdd.n648 37.0005
R3205 dvdd.n618 dvdd.n617 37.0005
R3206 dvdd.n617 dvdd.t30 37.0005
R3207 dvdd.n650 dvdd.n649 37.0005
R3208 dvdd.n649 dvdd.t19 37.0005
R3209 dvdd.n263 dvdd.n261 37.0005
R3210 dvdd.n597 dvdd.n262 33.2417
R3211 dvdd.n598 dvdd.n263 33.2417
R3212 dvdd.n564 dvdd.n553 31.2476
R3213 dvdd.n176 dvdd.n175 30.8338
R3214 dvdd.n175 dvdd.n154 30.8338
R3215 dvdd.n173 dvdd.n164 30.8338
R3216 dvdd.n173 dvdd.n154 30.8338
R3217 dvdd.n208 dvdd.n207 30.8338
R3218 dvdd.n208 dvdd.n154 30.8338
R3219 dvdd.n211 dvdd.n210 30.8338
R3220 dvdd.n210 dvdd.n154 30.8338
R3221 dvdd.n215 dvdd.n214 30.8338
R3222 dvdd.n214 dvdd.n154 30.8338
R3223 dvdd.n238 dvdd.n237 30.8338
R3224 dvdd.n237 dvdd.n135 30.8338
R3225 dvdd.n223 dvdd.n160 30.8338
R3226 dvdd.n160 dvdd.n154 30.8338
R3227 dvdd.n218 dvdd.n217 30.8338
R3228 dvdd.n217 dvdd.n134 30.8338
R3229 dvdd.n152 dvdd.n149 30.8338
R3230 dvdd.n152 dvdd.n134 30.8338
R3231 dvdd.n234 dvdd.n233 30.8338
R3232 dvdd.n234 dvdd.n135 30.8338
R3233 dvdd.n148 dvdd.n130 30.8338
R3234 dvdd.n135 dvdd.n130 30.8338
R3235 dvdd.n229 dvdd.n228 30.8338
R3236 dvdd.n228 dvdd.n134 30.8338
R3237 dvdd.n168 dvdd.n165 30.8338
R3238 dvdd.n168 dvdd.n134 30.8338
R3239 dvdd.n181 dvdd.n131 30.8338
R3240 dvdd.n135 dvdd.n131 30.8338
R3241 dvdd.n186 dvdd.n180 30.8338
R3242 dvdd.n180 dvdd.n135 30.8338
R3243 dvdd.n203 dvdd.n202 30.8338
R3244 dvdd.n202 dvdd.n134 30.8338
R3245 dvdd.n200 dvdd.n199 30.8338
R3246 dvdd.n200 dvdd.n134 30.8338
R3247 dvdd.n192 dvdd.n178 30.8338
R3248 dvdd.n192 dvdd.n135 30.8338
R3249 dvdd.n254 dvdd.n253 30.8338
R3250 dvdd.n255 dvdd.n254 30.8338
R3251 dvdd.n251 dvdd.n120 30.8338
R3252 dvdd.n255 dvdd.n120 30.8338
R3253 dvdd.n249 dvdd.n123 30.8338
R3254 dvdd.n255 dvdd.n123 30.8338
R3255 dvdd.n247 dvdd.n121 30.8338
R3256 dvdd.n255 dvdd.n121 30.8338
R3257 dvdd.n257 dvdd.n256 30.8338
R3258 dvdd.n256 dvdd.n255 30.8338
R3259 dvdd.n179 dvdd.n122 30.8338
R3260 dvdd.n255 dvdd.n122 30.8338
R3261 dvdd.n634 dvdd.n88 30.8338
R3262 dvdd.n634 dvdd.n70 30.8338
R3263 dvdd.n548 dvdd.n547 30.8338
R3264 dvdd.n547 dvdd.n56 30.8338
R3265 dvdd.n530 dvdd.n529 30.8338
R3266 dvdd.n529 dvdd.n55 30.8338
R3267 dvdd.n66 dvdd.n65 30.8338
R3268 dvdd.n65 dvdd.n56 30.8338
R3269 dvdd.n542 dvdd.n67 30.8338
R3270 dvdd.n542 dvdd.n56 30.8338
R3271 dvdd.n95 dvdd.n91 30.8338
R3272 dvdd.n95 dvdd.n55 30.8338
R3273 dvdd.n612 dvdd.n611 30.8338
R3274 dvdd.n611 dvdd.n97 30.8338
R3275 dvdd.n642 dvdd.n641 30.8338
R3276 dvdd.n642 dvdd.n79 30.8338
R3277 dvdd.n637 dvdd.n636 30.8338
R3278 dvdd.n636 dvdd.n70 30.8338
R3279 dvdd.n544 dvdd.n90 30.8338
R3280 dvdd.n544 dvdd.n56 30.8338
R3281 dvdd.n526 dvdd.n92 30.8338
R3282 dvdd.n526 dvdd.n55 30.8338
R3283 dvdd.n532 dvdd.n531 30.8338
R3284 dvdd.n532 dvdd.n97 30.8338
R3285 dvdd.n536 dvdd.n535 30.8338
R3286 dvdd.n535 dvdd.n97 30.8338
R3287 dvdd.n87 dvdd.n86 30.8338
R3288 dvdd.n86 dvdd.n79 30.8338
R3289 dvdd.n63 dvdd.n62 30.8338
R3290 dvdd.n62 dvdd.n55 30.8338
R3291 dvdd.n76 dvdd.n75 30.8338
R3292 dvdd.n75 dvdd.n70 30.8338
R3293 dvdd.n631 dvdd.n630 30.8338
R3294 dvdd.n631 dvdd.n70 30.8338
R3295 dvdd.n78 dvdd.n77 30.8338
R3296 dvdd.n79 dvdd.n78 30.8338
R3297 dvdd.n645 dvdd.n644 30.8338
R3298 dvdd.n644 dvdd.n79 30.8338
R3299 dvdd.n110 dvdd.n102 30.8338
R3300 dvdd.n110 dvdd.n97 30.8338
R3301 dvdd.n603 dvdd.n602 30.8338
R3302 dvdd.n602 dvdd.n105 30.8338
R3303 dvdd.n606 dvdd.n605 30.8338
R3304 dvdd.n606 dvdd.n105 30.8338
R3305 dvdd.n609 dvdd.n608 30.8338
R3306 dvdd.n608 dvdd.n105 30.8338
R3307 dvdd.n112 dvdd.n104 30.8338
R3308 dvdd.n105 dvdd.n104 30.8338
R3309 dvdd.n268 dvdd.n264 30.8338
R3310 dvdd.n525 dvdd.n524 30.8338
R3311 dvdd.n524 dvdd.n521 30.8338
R3312 dvdd.n583 dvdd.n273 30.8338
R3313 dvdd.n519 dvdd.n273 30.8338
R3314 dvdd.n591 dvdd.n267 30.8338
R3315 dvdd.n274 dvdd.n267 30.8338
R3316 dvdd.n564 dvdd.n554 30.8338
R3317 dvdd.n43 dvdd.n37 30.8338
R3318 dvdd.n39 dvdd.n36 30.8338
R3319 dvdd.n31 dvdd.n25 30.8338
R3320 dvdd.n27 dvdd.n24 30.8338
R3321 dvdd.n19 dvdd.n13 30.8338
R3322 dvdd.n15 dvdd.n12 30.8338
R3323 dvdd.n7 dvdd.n1 30.8338
R3324 dvdd.n3 dvdd.n0 30.8338
R3325 dvdd.n588 dvdd.n270 30.0837
R3326 dvdd.n587 dvdd.n586 25.7304
R3327 dvdd.n620 dvdd.n619 20.3196
R3328 dvdd.n620 dvdd.n51 20.3196
R3329 dvdd.n660 dvdd.n52 20.3196
R3330 dvdd.n652 dvdd.n52 20.3196
R3331 dvdd.n652 dvdd.n651 20.3196
R3332 dvdd.n586 dvdd.n585 20.2401
R3333 dvdd.n573 dvdd.n523 20.2401
R3334 dvdd.n661 dvdd.n51 17.1488
R3335 dvdd.n600 dvdd.n599 16.8187
R3336 dvdd.n596 dvdd.n595 16.8187
R3337 dvdd.n581 dvdd.n580 16.8187
R3338 dvdd.n585 dvdd.n584 16.8187
R3339 dvdd.n574 dvdd.n573 16.8187
R3340 dvdd.n570 dvdd.n569 16.8187
R3341 dvdd.n569 dvdd.t94 16.8187
R3342 dvdd.n567 dvdd.n566 16.8187
R3343 dvdd.n577 dvdd.n576 16.8187
R3344 dvdd.n576 dvdd.t119 16.8187
R3345 dvdd.n41 dvdd.n40 16.8187
R3346 dvdd.n45 dvdd.n44 16.8187
R3347 dvdd.n29 dvdd.n28 16.8187
R3348 dvdd.n33 dvdd.n32 16.8187
R3349 dvdd.n17 dvdd.n16 16.8187
R3350 dvdd.n21 dvdd.n20 16.8187
R3351 dvdd.n5 dvdd.n4 16.8187
R3352 dvdd.n9 dvdd.n8 16.8187
R3353 dvdd.n570 dvdd.n553 15.4969
R3354 dvdd.n573 dvdd.n572 14.3924
R3355 dvdd.n575 dvdd.n574 13.0425
R3356 dvdd.n584 dvdd.n272 13.0425
R3357 dvdd.n582 dvdd.n581 13.0425
R3358 dvdd.n568 dvdd.n567 13.0425
R3359 dvdd.n44 dvdd.n38 13.0425
R3360 dvdd.n42 dvdd.n41 13.0425
R3361 dvdd.n32 dvdd.n26 13.0425
R3362 dvdd.n30 dvdd.n29 13.0425
R3363 dvdd.n20 dvdd.n14 13.0425
R3364 dvdd.n18 dvdd.n17 13.0425
R3365 dvdd.n8 dvdd.n2 13.0425
R3366 dvdd.n6 dvdd.n5 13.0425
R3367 dvdd.n572 dvdd.n571 12.4107
R3368 dvdd.t89 dvdd.n357 11.9724
R3369 dvdd.n358 dvdd.t89 11.9724
R3370 dvdd.t0 dvdd.n379 11.9724
R3371 dvdd.n380 dvdd.t0 11.9724
R3372 dvdd.n270 dvdd.n264 11.3275
R3373 dvdd.n560 dvdd.n556 10.8829
R3374 dvdd.n557 dvdd.n518 10.8829
R3375 dvdd.n588 dvdd.n587 10.7538
R3376 dvdd.n585 dvdd.n271 10.6563
R3377 dvdd.n566 dvdd.n555 9.69349
R3378 dvdd.n558 dvdd.n557 9.61977
R3379 dvdd.n561 dvdd.n560 9.61977
R3380 dvdd.n523 dvdd.n271 9.58426
R3381 dvdd.n563 dvdd.n562 8.81002
R3382 dvdd.n559 dvdd.n275 8.81002
R3383 dvdd.n579 dvdd.n273 8.64212
R3384 dvdd.n267 dvdd.n265 8.64212
R3385 dvdd.n577 dvdd.n518 8.13999
R3386 dvdd.n523 dvdd.n273 8.08984
R3387 dvdd.n586 dvdd.n267 8.08984
R3388 dvdd.n241 dvdd.n240 7.4005
R3389 dvdd.t1 dvdd.n241 7.4005
R3390 dvdd.n219 dvdd.n140 7.4005
R3391 dvdd.t1 dvdd.n140 7.4005
R3392 dvdd.n231 dvdd.n139 7.4005
R3393 dvdd.t1 dvdd.n139 7.4005
R3394 dvdd.n242 dvdd.n133 7.4005
R3395 dvdd.n242 dvdd.t1 7.4005
R3396 dvdd.n166 dvdd.n138 7.4005
R3397 dvdd.t1 dvdd.n138 7.4005
R3398 dvdd.n187 dvdd.n137 7.4005
R3399 dvdd.t1 dvdd.n137 7.4005
R3400 dvdd.n197 dvdd.n136 7.4005
R3401 dvdd.t1 dvdd.n136 7.4005
R3402 dvdd.n593 dvdd.n592 7.4005
R3403 dvdd.n589 dvdd.n588 7.4005
R3404 dvdd.n601 dvdd.n260 7.31014
R3405 dvdd.n270 dvdd.n269 7.31014
R3406 dvdd.n253 dvdd.n252 6.58619
R3407 dvdd.n252 dvdd.n251 6.58619
R3408 dvdd.n251 dvdd.n250 6.58619
R3409 dvdd.n250 dvdd.n249 6.58619
R3410 dvdd.n249 dvdd.n248 6.58619
R3411 dvdd.n248 dvdd.n247 6.58619
R3412 dvdd.n247 dvdd.n116 6.58619
R3413 dvdd.n257 dvdd.n117 6.58619
R3414 dvdd.n179 dvdd.n117 6.58619
R3415 dvdd.n258 dvdd.n114 6.4005
R3416 dvdd.n578 dvdd.n577 6.36768
R3417 dvdd.n258 dvdd.n257 6.1653
R3418 dvdd.n486 dvdd.t50 5.91616
R3419 dvdd.t50 dvdd.n485 5.91616
R3420 dvdd.t14 dvdd.n503 5.91616
R3421 dvdd.n504 dvdd.t14 5.91616
R3422 dvdd.n512 dvdd.t25 5.91616
R3423 dvdd.t25 dvdd.n276 5.91616
R3424 dvdd.n458 dvdd.t43 5.91616
R3425 dvdd.t43 dvdd.n457 5.91616
R3426 dvdd.t56 dvdd.n481 5.91616
R3427 dvdd.n482 dvdd.t56 5.91616
R3428 dvdd.t65 dvdd.n440 5.91616
R3429 dvdd.n441 dvdd.t65 5.91616
R3430 dvdd.n590 dvdd.n589 5.51167
R3431 dvdd.n592 dvdd.n266 5.51167
R3432 dvdd.n485 dvdd.n484 5.13093
R3433 dvdd.n595 dvdd.n264 5.07987
R3434 dvdd.n423 dvdd.n422 4.88319
R3435 dvdd.n478 dvdd.n477 4.88319
R3436 dvdd.n49 dvdd.n48 4.88319
R3437 dvdd.n441 dvdd.n438 4.42713
R3438 dvdd.n483 dvdd.n482 4.42713
R3439 dvdd.n457 dvdd.n279 4.42713
R3440 dvdd.n458 dvdd.n277 4.42713
R3441 dvdd.n512 dvdd.n511 4.42713
R3442 dvdd.n504 dvdd.n282 4.42713
R3443 dvdd.n503 dvdd.n502 4.42713
R3444 dvdd.n485 dvdd.n297 4.42713
R3445 dvdd.n487 dvdd.n486 4.42713
R3446 dvdd.n481 dvdd.n480 4.38659
R3447 dvdd.n481 dvdd.n430 4.37758
R3448 dvdd.n440 dvdd.n432 4.37758
R3449 dvdd.n440 dvdd.n439 4.36463
R3450 dvdd.n442 dvdd.n441 4.36463
R3451 dvdd.n482 dvdd.n429 4.36463
R3452 dvdd.n457 dvdd.n456 4.36463
R3453 dvdd.n459 dvdd.n458 4.36463
R3454 dvdd.n513 dvdd.n512 4.36463
R3455 dvdd.n503 dvdd.n280 4.36463
R3456 dvdd.n486 dvdd.n296 4.36463
R3457 dvdd.n627 dvdd.n73 3.77601
R3458 dvdd.t44 dvdd.n73 3.77601
R3459 dvdd.n625 dvdd.n59 3.77601
R3460 dvdd.t26 dvdd.n59 3.77601
R3461 dvdd.n623 dvdd.n622 3.77601
R3462 dvdd.n622 dvdd.t15 3.77601
R3463 dvdd.n538 dvdd.n99 3.77601
R3464 dvdd.t15 dvdd.n99 3.77601
R3465 dvdd.n540 dvdd.n58 3.77601
R3466 dvdd.t26 dvdd.n58 3.77601
R3467 dvdd.n89 dvdd.n72 3.77601
R3468 dvdd.t44 dvdd.n72 3.77601
R3469 dvdd.n551 dvdd.n71 3.77601
R3470 dvdd.t44 dvdd.n71 3.77601
R3471 dvdd.n613 dvdd.n100 3.77601
R3472 dvdd.t15 dvdd.n100 3.77601
R3473 dvdd.n658 dvdd.n657 3.77601
R3474 dvdd.t26 dvdd.n658 3.77601
R3475 dvdd.n655 dvdd.n654 3.77601
R3476 dvdd.n654 dvdd.t44 3.77601
R3477 dvdd.n621 dvdd.n620 3.77601
R3478 dvdd.t15 dvdd.n621 3.77601
R3479 dvdd.n660 dvdd.n659 3.77601
R3480 dvdd.n659 dvdd.t26 3.77601
R3481 dvdd.n653 dvdd.n652 3.77601
R3482 dvdd.t44 dvdd.n653 3.77601
R3483 dvdd.n571 dvdd.n57 3.77601
R3484 dvdd.t26 dvdd.n57 3.77601
R3485 dvdd.n587 dvdd.n98 3.77601
R3486 dvdd.t15 dvdd.n98 3.77601
R3487 dvdd.t94 dvdd.n568 3.68792
R3488 dvdd.n582 dvdd.t106 3.68792
R3489 dvdd.t106 dvdd.n272 3.68792
R3490 dvdd.t119 dvdd.n575 3.68792
R3491 dvdd.n42 dvdd.t92 3.68792
R3492 dvdd.t92 dvdd.n38 3.68792
R3493 dvdd.n30 dvdd.t111 3.68792
R3494 dvdd.t111 dvdd.n26 3.68792
R3495 dvdd.n18 dvdd.t109 3.68792
R3496 dvdd.t109 dvdd.n14 3.68792
R3497 dvdd.n6 dvdd.t96 3.68792
R3498 dvdd.t96 dvdd.n2 3.68792
R3499 dvdd.n566 dvdd.n565 3.26067
R3500 dvdd.n598 dvdd.t99 3.25677
R3501 dvdd.t99 dvdd.n597 3.25677
R3502 dvdd.n661 dvdd.n660 3.17136
R3503 dvdd.n509 dvdd.n508 3.10376
R3504 dvdd.n516 dvdd.n515 3.04126
R3505 dvdd.n618 dvdd.n103 2.83329
R3506 dvdd.n619 dvdd.n618 2.83329
R3507 dvdd.n651 dvdd.n650 2.83329
R3508 dvdd.n506 dvdd.n505 2.74778
R3509 dvdd.n665 dvdd.n664 2.66096
R3510 dvdd.n420 dvdd.n419 2.42664
R3511 dvdd.n380 dvdd.n322 2.25322
R3512 dvdd.n379 dvdd.n378 2.25322
R3513 dvdd.n359 dvdd.n358 2.25322
R3514 dvdd.n357 dvdd.n354 2.25322
R3515 dvdd.n358 dvdd.n349 2.19072
R3516 dvdd.n357 dvdd.n356 2.19072
R3517 dvdd.n381 dvdd.n380 2.188
R3518 dvdd.n379 dvdd.n320 2.188
R3519 dvdd.n390 dvdd.n389 2.02496
R3520 dvdd.n571 dvdd.n570 1.98223
R3521 dvdd.t116 dvdd.n266 1.88064
R3522 dvdd.n590 dvdd.t116 1.88064
R3523 dvdd.n595 dvdd.n594 1.67669
R3524 dvdd.n555 dvdd.n518 1.554
R3525 dvdd.n505 dvdd.n504 1.37822
R3526 dvdd.n518 dvdd 1.3042
R3527 dvdd.n561 dvdd.t108 1.2275
R3528 dvdd.n558 dvdd.t108 1.2275
R3529 dvdd dvdd.n517 1.19558
R3530 dvdd.n508 dvdd.n276 1.08474
R3531 dvdd.n516 dvdd.n276 1.08474
R3532 dvdd.n517 dvdd.n516 0.996712
R3533 dvdd.n298 dvdd.n296 0.891804
R3534 dvdd.n418 dvdd.n417 0.860794
R3535 dvdd.n419 dvdd.n418 0.84943
R3536 dvdd.n484 dvdd.n483 0.791063
R3537 dvdd.n424 dvdd 0.751032
R3538 dvdd.n461 dvdd.n452 0.734196
R3539 dvdd.n329 dvdd.n328 0.734196
R3540 dvdd.n352 dvdd.n351 0.734196
R3541 dvdd.n47 dvdd.n46 0.639894
R3542 dvdd.n35 dvdd.n34 0.639894
R3543 dvdd.n23 dvdd.n22 0.639894
R3544 dvdd.n11 dvdd.n10 0.639894
R3545 dvdd dvdd.n667 0.62021
R3546 dvdd.n327 dvdd.n322 0.620065
R3547 dvdd.n378 dvdd.n377 0.620065
R3548 dvdd.n360 dvdd.n359 0.620065
R3549 dvdd.n354 dvdd.n353 0.620065
R3550 dvdd.n502 dvdd.n501 0.620065
R3551 dvdd.n297 dvdd.n290 0.620065
R3552 dvdd.n488 dvdd.n487 0.620065
R3553 dvdd.n426 dvdd.n425 0.603761
R3554 dvdd.n664 dvdd.n663 0.549667
R3555 dvdd.n476 dvdd.n475 0.478761
R3556 dvdd.n386 dvdd.n282 0.478761
R3557 dvdd.n421 dvdd.n293 0.478761
R3558 dvdd.n426 dvdd.n296 0.478761
R3559 dvdd.n425 dvdd.n421 0.474712
R3560 dvdd.n460 dvdd.n459 0.470609
R3561 dvdd.n438 dvdd.n429 0.470609
R3562 dvdd.n439 dvdd.n434 0.470609
R3563 dvdd.n443 dvdd.n442 0.470609
R3564 dvdd.n456 dvdd.n453 0.470609
R3565 dvdd.n513 dvdd.n279 0.470609
R3566 dvdd.n515 dvdd.n277 0.470609
R3567 dvdd.n511 dvdd.n280 0.470609
R3568 dvdd.n666 dvdd.n665 0.464907
R3569 dvdd.n667 dvdd.n666 0.464907
R3570 dvdd.n384 dvdd.n287 0.429848
R3571 dvdd.n445 dvdd.n443 0.429848
R3572 dvdd.n472 dvdd.n471 0.429848
R3573 dvdd.n449 dvdd.n447 0.429848
R3574 dvdd.n468 dvdd.n467 0.429848
R3575 dvdd.n453 dvdd.n451 0.429848
R3576 dvdd.n464 dvdd.n463 0.429848
R3577 dvdd.n331 dvdd.n330 0.429848
R3578 dvdd.n377 dvdd.n376 0.429848
R3579 dvdd.n335 dvdd.n333 0.429848
R3580 dvdd.n373 dvdd.n372 0.429848
R3581 dvdd.n339 dvdd.n337 0.429848
R3582 dvdd.n369 dvdd.n368 0.429848
R3583 dvdd.n343 dvdd.n341 0.429848
R3584 dvdd.n365 dvdd.n364 0.429848
R3585 dvdd.n350 dvdd.n345 0.429848
R3586 dvdd.n361 dvdd.n360 0.429848
R3587 dvdd.n304 dvdd.n302 0.429848
R3588 dvdd.n413 dvdd.n412 0.429848
R3589 dvdd.n308 dvdd.n306 0.429848
R3590 dvdd.n409 dvdd.n408 0.429848
R3591 dvdd.n312 dvdd.n310 0.429848
R3592 dvdd.n405 dvdd.n404 0.429848
R3593 dvdd.n317 dvdd.n314 0.429848
R3594 dvdd.n396 dvdd.n316 0.429848
R3595 dvdd.n394 dvdd.n393 0.429848
R3596 dvdd.n497 dvdd.n496 0.429848
R3597 dvdd.n501 dvdd.n500 0.429848
R3598 dvdd.n494 dvdd.n290 0.429848
R3599 dvdd.n492 dvdd.n491 0.429848
R3600 dvdd.n479 dvdd.n478 0.429489
R3601 dvdd.n258 dvdd.n116 0.42139
R3602 dvdd.n356 dvdd.n300 0.410826
R3603 dvdd.n349 dvdd.n302 0.410826
R3604 dvdd.n393 dvdd.n320 0.410826
R3605 dvdd.n382 dvdd.n381 0.410826
R3606 dvdd.n454 dvdd.n453 0.383652
R3607 dvdd.n460 dvdd.n454 0.383652
R3608 dvdd.n430 dvdd.n428 0.383652
R3609 dvdd.n483 dvdd.n428 0.383652
R3610 dvdd.n437 dvdd.n432 0.383652
R3611 dvdd.n438 dvdd.n437 0.383652
R3612 dvdd.n475 dvdd.n433 0.383652
R3613 dvdd.n472 dvdd.n433 0.383652
R3614 dvdd.n435 dvdd.n434 0.383652
R3615 dvdd.n443 dvdd.n435 0.383652
R3616 dvdd.n471 dvdd.n444 0.383652
R3617 dvdd.n468 dvdd.n444 0.383652
R3618 dvdd.n446 dvdd.n445 0.383652
R3619 dvdd.n447 dvdd.n446 0.383652
R3620 dvdd.n467 dvdd.n448 0.383652
R3621 dvdd.n464 dvdd.n448 0.383652
R3622 dvdd.n450 dvdd.n449 0.383652
R3623 dvdd.n451 dvdd.n450 0.383652
R3624 dvdd.n463 dvdd.n452 0.383652
R3625 dvdd.n279 dvdd.n278 0.383652
R3626 dvdd.n278 dvdd.n277 0.383652
R3627 dvdd.n511 dvdd.n510 0.383652
R3628 dvdd.n510 dvdd.n509 0.383652
R3629 dvdd.n313 dvdd.n312 0.383652
R3630 dvdd.n314 dvdd.n313 0.383652
R3631 dvdd.n330 dvdd.n329 0.383652
R3632 dvdd.n377 dvdd.n324 0.383652
R3633 dvdd.n327 dvdd.n324 0.383652
R3634 dvdd.n378 dvdd.n323 0.383652
R3635 dvdd.n323 dvdd.n322 0.383652
R3636 dvdd.n373 dvdd.n326 0.383652
R3637 dvdd.n376 dvdd.n326 0.383652
R3638 dvdd.n333 dvdd.n332 0.383652
R3639 dvdd.n332 dvdd.n331 0.383652
R3640 dvdd.n369 dvdd.n334 0.383652
R3641 dvdd.n372 dvdd.n334 0.383652
R3642 dvdd.n337 dvdd.n336 0.383652
R3643 dvdd.n336 dvdd.n335 0.383652
R3644 dvdd.n365 dvdd.n338 0.383652
R3645 dvdd.n368 dvdd.n338 0.383652
R3646 dvdd.n341 dvdd.n340 0.383652
R3647 dvdd.n340 dvdd.n339 0.383652
R3648 dvdd.n361 dvdd.n342 0.383652
R3649 dvdd.n364 dvdd.n342 0.383652
R3650 dvdd.n345 dvdd.n344 0.383652
R3651 dvdd.n344 dvdd.n343 0.383652
R3652 dvdd.n353 dvdd.n346 0.383652
R3653 dvdd.n360 dvdd.n346 0.383652
R3654 dvdd.n354 dvdd.n348 0.383652
R3655 dvdd.n359 dvdd.n348 0.383652
R3656 dvdd.n351 dvdd.n350 0.383652
R3657 dvdd.n416 dvdd.n299 0.383652
R3658 dvdd.n413 dvdd.n299 0.383652
R3659 dvdd.n301 dvdd.n300 0.383652
R3660 dvdd.n302 dvdd.n301 0.383652
R3661 dvdd.n412 dvdd.n303 0.383652
R3662 dvdd.n409 dvdd.n303 0.383652
R3663 dvdd.n305 dvdd.n304 0.383652
R3664 dvdd.n306 dvdd.n305 0.383652
R3665 dvdd.n408 dvdd.n307 0.383652
R3666 dvdd.n405 dvdd.n307 0.383652
R3667 dvdd.n309 dvdd.n308 0.383652
R3668 dvdd.n310 dvdd.n309 0.383652
R3669 dvdd.n404 dvdd.n311 0.383652
R3670 dvdd.n400 dvdd.n311 0.383652
R3671 dvdd.n318 dvdd.n317 0.383652
R3672 dvdd.n394 dvdd.n318 0.383652
R3673 dvdd.n400 dvdd.n397 0.383652
R3674 dvdd.n397 dvdd.n396 0.383652
R3675 dvdd.n393 dvdd.n319 0.383652
R3676 dvdd.n382 dvdd.n319 0.383652
R3677 dvdd.n383 dvdd.n316 0.383652
R3678 dvdd.n390 dvdd.n383 0.383652
R3679 dvdd.n385 dvdd.n384 0.383652
R3680 dvdd.n389 dvdd.n385 0.383652
R3681 dvdd.n501 dvdd.n284 0.383652
R3682 dvdd.n387 dvdd.n284 0.383652
R3683 dvdd.n502 dvdd.n283 0.383652
R3684 dvdd.n283 dvdd.n282 0.383652
R3685 dvdd.n497 dvdd.n286 0.383652
R3686 dvdd.n500 dvdd.n286 0.383652
R3687 dvdd.n492 dvdd.n291 0.383652
R3688 dvdd.n399 dvdd.n291 0.383652
R3689 dvdd.n399 dvdd.n398 0.383652
R3690 dvdd.n398 dvdd.n287 0.383652
R3691 dvdd.n495 dvdd.n494 0.383652
R3692 dvdd.n496 dvdd.n495 0.383652
R3693 dvdd.n293 dvdd.n292 0.383652
R3694 dvdd.n491 dvdd.n292 0.383652
R3695 dvdd.n487 dvdd.n295 0.383652
R3696 dvdd.n297 dvdd.n295 0.383652
R3697 dvdd.n488 dvdd.n294 0.383652
R3698 dvdd.n294 dvdd.n290 0.383652
R3699 dvdd.n420 dvdd.n416 0.373755
R3700 dvdd.n484 dvdd.n427 0.373227
R3701 dvdd.n400 dvdd.n399 0.373
R3702 dvdd.n461 dvdd.n460 0.351043
R3703 dvdd.n474 dvdd.n434 0.351043
R3704 dvdd.n475 dvdd.n474 0.351043
R3705 dvdd.n473 dvdd.n443 0.351043
R3706 dvdd.n473 dvdd.n472 0.351043
R3707 dvdd.n470 dvdd.n445 0.351043
R3708 dvdd.n471 dvdd.n470 0.351043
R3709 dvdd.n469 dvdd.n447 0.351043
R3710 dvdd.n469 dvdd.n468 0.351043
R3711 dvdd.n466 dvdd.n449 0.351043
R3712 dvdd.n467 dvdd.n466 0.351043
R3713 dvdd.n465 dvdd.n451 0.351043
R3714 dvdd.n465 dvdd.n464 0.351043
R3715 dvdd.n462 dvdd.n453 0.351043
R3716 dvdd.n463 dvdd.n462 0.351043
R3717 dvdd.n328 dvdd.n327 0.351043
R3718 dvdd.n330 dvdd.n325 0.351043
R3719 dvdd.n377 dvdd.n325 0.351043
R3720 dvdd.n375 dvdd.n331 0.351043
R3721 dvdd.n376 dvdd.n375 0.351043
R3722 dvdd.n374 dvdd.n333 0.351043
R3723 dvdd.n374 dvdd.n373 0.351043
R3724 dvdd.n371 dvdd.n335 0.351043
R3725 dvdd.n372 dvdd.n371 0.351043
R3726 dvdd.n370 dvdd.n337 0.351043
R3727 dvdd.n370 dvdd.n369 0.351043
R3728 dvdd.n367 dvdd.n339 0.351043
R3729 dvdd.n368 dvdd.n367 0.351043
R3730 dvdd.n366 dvdd.n341 0.351043
R3731 dvdd.n366 dvdd.n365 0.351043
R3732 dvdd.n363 dvdd.n343 0.351043
R3733 dvdd.n364 dvdd.n363 0.351043
R3734 dvdd.n362 dvdd.n345 0.351043
R3735 dvdd.n362 dvdd.n361 0.351043
R3736 dvdd.n350 dvdd.n347 0.351043
R3737 dvdd.n360 dvdd.n347 0.351043
R3738 dvdd.n353 dvdd.n352 0.351043
R3739 dvdd.n415 dvdd.n300 0.351043
R3740 dvdd.n416 dvdd.n415 0.351043
R3741 dvdd.n414 dvdd.n302 0.351043
R3742 dvdd.n414 dvdd.n413 0.351043
R3743 dvdd.n411 dvdd.n304 0.351043
R3744 dvdd.n412 dvdd.n411 0.351043
R3745 dvdd.n410 dvdd.n306 0.351043
R3746 dvdd.n410 dvdd.n409 0.351043
R3747 dvdd.n407 dvdd.n308 0.351043
R3748 dvdd.n408 dvdd.n407 0.351043
R3749 dvdd.n406 dvdd.n310 0.351043
R3750 dvdd.n406 dvdd.n405 0.351043
R3751 dvdd.n403 dvdd.n312 0.351043
R3752 dvdd.n404 dvdd.n403 0.351043
R3753 dvdd.n402 dvdd.n314 0.351043
R3754 dvdd.n317 dvdd.n315 0.351043
R3755 dvdd.n395 dvdd.n394 0.351043
R3756 dvdd.n396 dvdd.n395 0.351043
R3757 dvdd.n393 dvdd.n392 0.351043
R3758 dvdd.n392 dvdd.n316 0.351043
R3759 dvdd.n391 dvdd.n382 0.351043
R3760 dvdd.n391 dvdd.n390 0.351043
R3761 dvdd.n389 dvdd.n388 0.351043
R3762 dvdd.n388 dvdd.n387 0.351043
R3763 dvdd.n384 dvdd.n285 0.351043
R3764 dvdd.n501 dvdd.n285 0.351043
R3765 dvdd.n498 dvdd.n497 0.351043
R3766 dvdd.n499 dvdd.n287 0.351043
R3767 dvdd.n500 dvdd.n499 0.351043
R3768 dvdd.n496 dvdd.n289 0.351043
R3769 dvdd.n493 dvdd.n492 0.351043
R3770 dvdd.n494 dvdd.n493 0.351043
R3771 dvdd.n491 dvdd.n490 0.351043
R3772 dvdd.n490 dvdd.n290 0.351043
R3773 dvdd.n489 dvdd.n293 0.351043
R3774 dvdd.n489 dvdd.n488 0.351043
R3775 dvdd.n507 dvdd.n506 0.307565
R3776 dvdd.n402 dvdd.n401 0.288543
R3777 dvdd.n401 dvdd.n315 0.288543
R3778 dvdd.n498 dvdd.n288 0.288543
R3779 dvdd.n289 dvdd.n288 0.288543
R3780 dvdd.n439 dvdd.n436 0.263321
R3781 dvdd.n442 dvdd.n436 0.263321
R3782 dvdd.n431 dvdd.n429 0.263321
R3783 dvdd.n456 dvdd.n455 0.263321
R3784 dvdd.n459 dvdd.n455 0.263321
R3785 dvdd.n514 dvdd.n513 0.263321
R3786 dvdd.n515 dvdd.n514 0.263321
R3787 dvdd.n281 dvdd.n280 0.263321
R3788 dvdd.n506 dvdd.n281 0.263321
R3789 dvdd.n480 dvdd.n431 0.226462
R3790 dvdd.n356 dvdd.n355 0.2055
R3791 dvdd.n355 dvdd.n349 0.2055
R3792 dvdd.n321 dvdd.n320 0.20347
R3793 dvdd.n381 dvdd.n321 0.20347
R3794 dvdd.n252 dvdd.n103 0.198679
R3795 dvdd.n663 dvdd 0.177824
R3796 dvdd.n663 dvdd.n49 0.170597
R3797 dvdd.n509 dvdd.n507 0.163543
R3798 dvdd.n665 dvdd 0.155803
R3799 dvdd.n666 dvdd 0.155803
R3800 dvdd.n667 dvdd 0.155803
R3801 dvdd.n387 dvdd.n386 0.141804
R3802 dvdd.n484 dvdd.n298 0.1255
R3803 dvdd.n479 dvdd.n432 0.0646892
R3804 dvdd.n478 dvdd.n476 0.0616026
R3805 dvdd.n421 dvdd.n420 0.0612215
R3806 dvdd.n430 dvdd.n50 0.0579324
R3807 dvdd.n480 dvdd.n479 0.0556802
R3808 dvdd.n427 dvdd.n50 0.0556802
R3809 dvdd.n46 dvdd.n45 0.0556724
R3810 dvdd.n34 dvdd.n33 0.0556724
R3811 dvdd.n22 dvdd.n21 0.0556724
R3812 dvdd.n10 dvdd.n9 0.0556724
R3813 dvdd.n662 dvdd.n50 0.0414555
R3814 dvdd dvdd.n47 0.0390101
R3815 dvdd dvdd.n35 0.0390101
R3816 dvdd dvdd.n23 0.0390101
R3817 dvdd dvdd.n11 0.0390101
R3818 dvdd.n269 dvdd.n260 0.0329873
R3819 dvdd.n662 dvdd.n661 0.0196358
R3820 dvdd.n476 dvdd 0.0171413
R3821 dvdd.n663 dvdd.n662 0.0165004
R3822 dvdd.n427 dvdd.n426 0.0162658
R3823 dvdd.n479 dvdd.n49 0.0139654
R3824 dvdd.n401 dvdd.n400 0.012
R3825 dvdd.n399 dvdd.n288 0.012
R3826 dvdd.n664 dvdd 0.0109536
R3827 dvdd.n423 dvdd.n50 0.00386852
R3828 dvdd.n425 dvdd.n424 0.00189736
R3829 dvdd.n424 dvdd.n423 0.000668426
R3830 comp_hyst_0.net3.t0 comp_hyst_0.net3.t1 242.977
R3831 comp_hyst_0.net3.t0 comp_hyst_0.net3.t3 242.409
R3832 comp_hyst_0.net3.t0 comp_hyst_0.net3.t2 230.071
R3833 level_shifter_3.in_b.t0 level_shifter_3.in_b.t1 229.644
R3834 level_shifter_3.in_b.t2 level_shifter_3.in_b.t0 27.1253
R3835 multiplexer_0.vtrip_3.n0 multiplexer_0.vtrip_3.t1 227.385
R3836 multiplexer_0.trans_gate_m_33.ena_b multiplexer_0.vtrip_3.t4 97.296
R3837 multiplexer_0.vtrip_3.n0 multiplexer_0.vtrip_3.t0 41.2565
R3838 multiplexer_0.vtrip_3.n0 multiplexer_0.trans_gate_m_33.ena_b 27.5547
R3839 multiplexer_0.trans_gate_m_33.ena_b multiplexer_0.vtrip_3.t5 18.5516
R3840 multiplexer_0.trans_gate_m_33.ena_b multiplexer_0.vtrip_3.t3 18.1873
R3841 multiplexer_0.vtrip_3.n0 multiplexer_0.vtrip_3.t2 16.8956
R3842 multiplexer_0.in_0110.n0 multiplexer_0.in_0110.t2 228.216
R3843 multiplexer_0.in_0110.n0 multiplexer_0.in_0110.t1 83.695
R3844 multiplexer_0.in_0110.n4 multiplexer_0.in_0110.t0 10.5295
R3845 multiplexer_0.in_0110.n4 multiplexer_0.in_0110.t3 10.5285
R3846 multiplexer_0.in_0110 multiplexer_0.in_0110.n3 4.51461
R3847 multiplexer_0.in_0110.n2 multiplexer_0.in_0110.n1 4.34635
R3848 multiplexer_0.in_0110.n1 multiplexer_0.in_0110.n0 1.5005
R3849 multiplexer_0.in_0110 multiplexer_0.in_0110.n4 0.872792
R3850 multiplexer_0.in_0110.n3 multiplexer_0.in_0110 0.177654
R3851 multiplexer_0.in_0110.n1 multiplexer_0.in_0110 0.104667
R3852 multiplexer_0.in_0110.n2 multiplexer_0.in_0110 0.0064902
R3853 multiplexer_0.in_0110.n3 multiplexer_0.in_0110.n2 0.00411538
R3854 level_shifter_2.out multiplexer_0.vtrip_2.t0 227.385
R3855 multiplexer_0.trans_gate_m_20.ena_b multiplexer_0.vtrip_2.t1 97.296
R3856 multiplexer_0.trans_gate_m_20.ena_b multiplexer_0.vtrip_2.n0 20.952
R3857 level_shifter_2.out multiplexer_0.trans_gate_m_20.ena_b 20.7215
R3858 multiplexer_0.trans_gate_m_20.ena_b multiplexer_0.vtrip_2.t3 18.5516
R3859 multiplexer_0.trans_gate_m_20.ena_b multiplexer_0.vtrip_2.t6 18.1873
R3860 level_shifter_2.out multiplexer_0.vtrip_2.t5 16.8956
R3861 multiplexer_0.vtrip_2.n0 multiplexer_0.vtrip_2.t2 16.8731
R3862 multiplexer_0.vtrip_2.n0 multiplexer_0.vtrip_2.t4 16.5088
R3863 multiplexer_0.in_1100.n0 multiplexer_0.in_1100.t1 228.216
R3864 multiplexer_0.in_1100.n0 multiplexer_0.in_1100.t2 83.695
R3865 multiplexer_0.in_1100.n3 multiplexer_0.in_1100.t3 10.5739
R3866 multiplexer_0.in_1100.n3 multiplexer_0.in_1100.t0 10.5739
R3867 multiplexer_0.in_1100 multiplexer_0.in_1100.n3 2.20538
R3868 multiplexer_0.in_1100 multiplexer_0.in_1100.n0 1.60467
R3869 multiplexer_0.in_1100 multiplexer_0.in_1100.n2 0.9755
R3870 multiplexer_0.in_1100.n2 multiplexer_0.in_1100 0.471654
R3871 multiplexer_0.in_1100.n1 multiplexer_0.in_1100 0.414042
R3872 multiplexer_0.in_1100.n1 multiplexer_0.in_1100 0.0140417
R3873 multiplexer_0.in_1100.n2 multiplexer_0.in_1100.n1 0.0101154
R3874 multiplexer_0.in_1101.n0 multiplexer_0.in_1101.t0 228.216
R3875 multiplexer_0.in_1101.n0 multiplexer_0.in_1101.t1 83.695
R3876 multiplexer_0.in_1101.n3 multiplexer_0.in_1101.t2 10.5295
R3877 multiplexer_0.in_1101.n3 multiplexer_0.in_1101.t3 10.5285
R3878 multiplexer_0.in_1101 multiplexer_0.in_1101.n2 3.98817
R3879 multiplexer_0.in_1101 multiplexer_0.in_1101.n0 1.60467
R3880 multiplexer_0.in_1101 multiplexer_0.in_1101.n3 0.872792
R3881 multiplexer_0.in_1101.n2 multiplexer_0.in_1101 0.471654
R3882 multiplexer_0.in_1101.n1 multiplexer_0.in_1101 0.414042
R3883 multiplexer_0.in_1101.n1 multiplexer_0.in_1101 0.0140417
R3884 multiplexer_0.in_1101.n2 multiplexer_0.in_1101.n1 0.0101154
R3885 vtrip[0].n2 vtrip[0].t2 99.4021
R3886 vtrip[0].n0 vtrip[0].t1 23.1698
R3887 vtrip[0].n1 vtrip[0].t3 17.7681
R3888 vtrip[0].n0 vtrip[0].t0 17.7475
R3889 vtrip[0].n2 vtrip[0] 5.62823
R3890 vtrip[0].n3 vtrip[0].n2 1.7055
R3891 vtrip[0].n1 vtrip[0].n0 0.572059
R3892 vtrip[0].n3 vtrip[0].n1 0.1139
R3893 vtrip[0] vtrip[0].n3 0.0378665
R3894 level_shifter_0.in_b.t1 level_shifter_0.in_b.t0 229.644
R3895 level_shifter_0.in_b.t2 level_shifter_0.in_b.t1 27.1253
R3896 multiplexer_0.trans_gate_m_32.in.t0 multiplexer_0.trans_gate_m_32.in.t2 228.216
R3897 multiplexer_0.trans_gate_m_32.in.t0 multiplexer_0.trans_gate_m_32.in.t4 228.216
R3898 multiplexer_0.trans_gate_m_32.in.t0 multiplexer_0.trans_gate_m_32.in.t1 228.216
R3899 multiplexer_0.trans_gate_m_32.in.t0 multiplexer_0.trans_gate_m_32.in.t3 93.748
R3900 multiplexer_0.trans_gate_m_37.out.t3 multiplexer_0.trans_gate_m_37.out.t2 228.216
R3901 multiplexer_0.trans_gate_m_37.out.t3 multiplexer_0.trans_gate_m_37.out.t5 228.216
R3902 multiplexer_0.trans_gate_m_37.out.t3 multiplexer_0.trans_gate_m_37.out.t1 228.216
R3903 multiplexer_0.trans_gate_m_37.out.t3 multiplexer_0.trans_gate_m_37.out.t4 94.7343
R3904 multiplexer_0.trans_gate_m_37.out.t3 multiplexer_0.trans_gate_m_37.out.t0 83.695
R3905 avdd.n84 avdd.n78 1446.62
R3906 avdd.n81 avdd.n80 1446.62
R3907 avdd.n73 avdd.n67 1446.62
R3908 avdd.n70 avdd.n69 1446.62
R3909 avdd.n62 avdd.n56 1446.62
R3910 avdd.n59 avdd.n58 1446.62
R3911 avdd.n51 avdd.n45 1446.62
R3912 avdd.n48 avdd.n47 1446.62
R3913 avdd.n40 avdd.n34 1446.62
R3914 avdd.n37 avdd.n36 1446.62
R3915 avdd.n29 avdd.n23 1446.62
R3916 avdd.n26 avdd.n25 1446.62
R3917 avdd.n18 avdd.n12 1446.62
R3918 avdd.n15 avdd.n14 1446.62
R3919 avdd.n7 avdd.n1 1446.62
R3920 avdd.n4 avdd.n3 1446.62
R3921 avdd.n172 avdd.n166 1446.62
R3922 avdd.n169 avdd.n168 1446.62
R3923 avdd.n161 avdd.n155 1446.62
R3924 avdd.n158 avdd.n157 1446.62
R3925 avdd.n150 avdd.n144 1446.62
R3926 avdd.n147 avdd.n146 1446.62
R3927 avdd.n139 avdd.n133 1446.62
R3928 avdd.n136 avdd.n135 1446.62
R3929 avdd.n128 avdd.n122 1446.62
R3930 avdd.n125 avdd.n124 1446.62
R3931 avdd.n117 avdd.n111 1446.62
R3932 avdd.n114 avdd.n113 1446.62
R3933 avdd.n106 avdd.n100 1446.62
R3934 avdd.n103 avdd.n102 1446.62
R3935 avdd.n95 avdd.n89 1446.62
R3936 avdd.n92 avdd.n91 1446.62
R3937 avdd.n260 avdd.n254 1446.62
R3938 avdd.n257 avdd.n256 1446.62
R3939 avdd.n249 avdd.n243 1446.62
R3940 avdd.n246 avdd.n245 1446.62
R3941 avdd.n238 avdd.n232 1446.62
R3942 avdd.n235 avdd.n234 1446.62
R3943 avdd.n227 avdd.n221 1446.62
R3944 avdd.n224 avdd.n223 1446.62
R3945 avdd.n216 avdd.n210 1446.62
R3946 avdd.n213 avdd.n212 1446.62
R3947 avdd.n205 avdd.n199 1446.62
R3948 avdd.n202 avdd.n201 1446.62
R3949 avdd.n194 avdd.n188 1446.62
R3950 avdd.n191 avdd.n190 1446.62
R3951 avdd.n183 avdd.n177 1446.62
R3952 avdd.n180 avdd.n179 1446.62
R3953 avdd.n304 avdd.n298 1446.62
R3954 avdd.n301 avdd.n300 1446.62
R3955 avdd.n293 avdd.n287 1446.62
R3956 avdd.n290 avdd.n289 1446.62
R3957 avdd.n282 avdd.n276 1446.62
R3958 avdd.n279 avdd.n278 1446.62
R3959 avdd.n271 avdd.n265 1446.62
R3960 avdd.n268 avdd.n267 1446.62
R3961 avdd.n326 avdd.n319 1446.62
R3962 avdd.n326 avdd.n317 1446.62
R3963 avdd.n327 avdd.n311 1446.62
R3964 avdd.n327 avdd.n312 1446.62
R3965 avdd.n349 avdd.n342 1446.62
R3966 avdd.n349 avdd.n340 1446.62
R3967 avdd.n350 avdd.n334 1446.62
R3968 avdd.n350 avdd.n335 1446.62
R3969 avdd.n373 avdd.n366 1446.62
R3970 avdd.n373 avdd.n364 1446.62
R3971 avdd.n374 avdd.n358 1446.62
R3972 avdd.n374 avdd.n359 1446.62
R3973 avdd.n397 avdd.n390 1446.62
R3974 avdd.n397 avdd.n388 1446.62
R3975 avdd.n398 avdd.n382 1446.62
R3976 avdd.n398 avdd.n383 1446.62
R3977 avdd.n316 avdd.n314 910.034
R3978 avdd.n318 avdd.n314 910.034
R3979 avdd.n339 avdd.n337 910.034
R3980 avdd.n341 avdd.n337 910.034
R3981 avdd.n363 avdd.n361 910.034
R3982 avdd.n365 avdd.n361 910.034
R3983 avdd.n387 avdd.n385 910.034
R3984 avdd.n389 avdd.n385 910.034
R3985 avdd.n319 avdd.n318 536.587
R3986 avdd.n316 avdd.n311 536.587
R3987 avdd.n317 avdd.n316 536.587
R3988 avdd.n318 avdd.n312 536.587
R3989 avdd.n342 avdd.n341 536.587
R3990 avdd.n339 avdd.n334 536.587
R3991 avdd.n340 avdd.n339 536.587
R3992 avdd.n341 avdd.n335 536.587
R3993 avdd.n366 avdd.n365 536.587
R3994 avdd.n363 avdd.n358 536.587
R3995 avdd.n364 avdd.n363 536.587
R3996 avdd.n365 avdd.n359 536.587
R3997 avdd.n390 avdd.n389 536.587
R3998 avdd.n387 avdd.n382 536.587
R3999 avdd.n388 avdd.n387 536.587
R4000 avdd.n389 avdd.n383 536.587
R4001 avdd.n82 avdd.n78 410.803
R4002 avdd.n83 avdd.n80 410.803
R4003 avdd.n71 avdd.n67 410.803
R4004 avdd.n72 avdd.n69 410.803
R4005 avdd.n60 avdd.n56 410.803
R4006 avdd.n61 avdd.n58 410.803
R4007 avdd.n49 avdd.n45 410.803
R4008 avdd.n50 avdd.n47 410.803
R4009 avdd.n38 avdd.n34 410.803
R4010 avdd.n39 avdd.n36 410.803
R4011 avdd.n27 avdd.n23 410.803
R4012 avdd.n28 avdd.n25 410.803
R4013 avdd.n16 avdd.n12 410.803
R4014 avdd.n17 avdd.n14 410.803
R4015 avdd.n5 avdd.n1 410.803
R4016 avdd.n6 avdd.n3 410.803
R4017 avdd.n170 avdd.n166 410.803
R4018 avdd.n171 avdd.n168 410.803
R4019 avdd.n159 avdd.n155 410.803
R4020 avdd.n160 avdd.n157 410.803
R4021 avdd.n148 avdd.n144 410.803
R4022 avdd.n149 avdd.n146 410.803
R4023 avdd.n137 avdd.n133 410.803
R4024 avdd.n138 avdd.n135 410.803
R4025 avdd.n126 avdd.n122 410.803
R4026 avdd.n127 avdd.n124 410.803
R4027 avdd.n115 avdd.n111 410.803
R4028 avdd.n116 avdd.n113 410.803
R4029 avdd.n104 avdd.n100 410.803
R4030 avdd.n105 avdd.n102 410.803
R4031 avdd.n93 avdd.n89 410.803
R4032 avdd.n94 avdd.n91 410.803
R4033 avdd.n258 avdd.n254 410.803
R4034 avdd.n259 avdd.n256 410.803
R4035 avdd.n247 avdd.n243 410.803
R4036 avdd.n248 avdd.n245 410.803
R4037 avdd.n236 avdd.n232 410.803
R4038 avdd.n237 avdd.n234 410.803
R4039 avdd.n225 avdd.n221 410.803
R4040 avdd.n226 avdd.n223 410.803
R4041 avdd.n214 avdd.n210 410.803
R4042 avdd.n215 avdd.n212 410.803
R4043 avdd.n203 avdd.n199 410.803
R4044 avdd.n204 avdd.n201 410.803
R4045 avdd.n192 avdd.n188 410.803
R4046 avdd.n193 avdd.n190 410.803
R4047 avdd.n181 avdd.n177 410.803
R4048 avdd.n182 avdd.n179 410.803
R4049 avdd.n302 avdd.n298 410.803
R4050 avdd.n303 avdd.n300 410.803
R4051 avdd.n291 avdd.n287 410.803
R4052 avdd.n292 avdd.n289 410.803
R4053 avdd.n280 avdd.n276 410.803
R4054 avdd.n281 avdd.n278 410.803
R4055 avdd.n269 avdd.n265 410.803
R4056 avdd.n270 avdd.n267 410.803
R4057 avdd.t16 avdd.n313 314.628
R4058 avdd.t16 avdd.n315 314.628
R4059 avdd.t5 avdd.n336 314.628
R4060 avdd.t5 avdd.n338 314.628
R4061 avdd.t28 avdd.n360 314.628
R4062 avdd.t28 avdd.n362 314.628
R4063 avdd.t21 avdd.n384 314.628
R4064 avdd.t21 avdd.n386 314.628
R4065 avdd.n85 avdd.n79 281.601
R4066 avdd.n74 avdd.n68 281.601
R4067 avdd.n63 avdd.n57 281.601
R4068 avdd.n52 avdd.n46 281.601
R4069 avdd.n41 avdd.n35 281.601
R4070 avdd.n30 avdd.n24 281.601
R4071 avdd.n19 avdd.n13 281.601
R4072 avdd.n8 avdd.n2 281.601
R4073 avdd.n173 avdd.n167 281.601
R4074 avdd.n162 avdd.n156 281.601
R4075 avdd.n151 avdd.n145 281.601
R4076 avdd.n140 avdd.n134 281.601
R4077 avdd.n129 avdd.n123 281.601
R4078 avdd.n118 avdd.n112 281.601
R4079 avdd.n107 avdd.n101 281.601
R4080 avdd.n96 avdd.n90 281.601
R4081 avdd.n261 avdd.n255 281.601
R4082 avdd.n250 avdd.n244 281.601
R4083 avdd.n239 avdd.n233 281.601
R4084 avdd.n228 avdd.n222 281.601
R4085 avdd.n217 avdd.n211 281.601
R4086 avdd.n206 avdd.n200 281.601
R4087 avdd.n195 avdd.n189 281.601
R4088 avdd.n184 avdd.n178 281.601
R4089 avdd.n305 avdd.n299 281.601
R4090 avdd.n294 avdd.n288 281.601
R4091 avdd.n283 avdd.n277 281.601
R4092 avdd.n272 avdd.n266 281.601
R4093 avdd.n308 avdd.t27 227.845
R4094 avdd.n331 avdd.t6 227.845
R4095 avdd.n355 avdd.t37 227.845
R4096 avdd.n379 avdd.t25 227.845
R4097 avdd.n308 avdd.t17 227.345
R4098 avdd.n331 avdd.t10 227.345
R4099 avdd.n355 avdd.t29 227.345
R4100 avdd.n379 avdd.t22 227.345
R4101 avdd.n79 avdd.n77 217.418
R4102 avdd.n68 avdd.n66 217.418
R4103 avdd.n57 avdd.n55 217.418
R4104 avdd.n46 avdd.n44 217.418
R4105 avdd.n35 avdd.n33 217.418
R4106 avdd.n24 avdd.n22 217.418
R4107 avdd.n13 avdd.n11 217.418
R4108 avdd.n2 avdd.n0 217.418
R4109 avdd.n167 avdd.n165 217.418
R4110 avdd.n156 avdd.n154 217.418
R4111 avdd.n145 avdd.n143 217.418
R4112 avdd.n134 avdd.n132 217.418
R4113 avdd.n123 avdd.n121 217.418
R4114 avdd.n112 avdd.n110 217.418
R4115 avdd.n101 avdd.n99 217.418
R4116 avdd.n90 avdd.n88 217.418
R4117 avdd.n255 avdd.n253 217.418
R4118 avdd.n244 avdd.n242 217.418
R4119 avdd.n233 avdd.n231 217.418
R4120 avdd.n222 avdd.n220 217.418
R4121 avdd.n211 avdd.n209 217.418
R4122 avdd.n200 avdd.n198 217.418
R4123 avdd.n189 avdd.n187 217.418
R4124 avdd.n178 avdd.n176 217.418
R4125 avdd.n299 avdd.n297 217.418
R4126 avdd.n288 avdd.n286 217.418
R4127 avdd.n277 avdd.n275 217.418
R4128 avdd.n266 avdd.n264 217.418
R4129 avdd.n86 avdd.n85 205.571
R4130 avdd.n75 avdd.n74 205.571
R4131 avdd.n64 avdd.n63 205.571
R4132 avdd.n53 avdd.n52 205.571
R4133 avdd.n42 avdd.n41 205.571
R4134 avdd.n31 avdd.n30 205.571
R4135 avdd.n20 avdd.n19 205.571
R4136 avdd.n9 avdd.n8 205.571
R4137 avdd.n174 avdd.n173 205.571
R4138 avdd.n163 avdd.n162 205.571
R4139 avdd.n152 avdd.n151 205.571
R4140 avdd.n141 avdd.n140 205.571
R4141 avdd.n130 avdd.n129 205.571
R4142 avdd.n119 avdd.n118 205.571
R4143 avdd.n108 avdd.n107 205.571
R4144 avdd.n97 avdd.n96 205.571
R4145 avdd.n262 avdd.n261 205.571
R4146 avdd.n251 avdd.n250 205.571
R4147 avdd.n240 avdd.n239 205.571
R4148 avdd.n229 avdd.n228 205.571
R4149 avdd.n218 avdd.n217 205.571
R4150 avdd.n207 avdd.n206 205.571
R4151 avdd.n196 avdd.n195 205.571
R4152 avdd.n185 avdd.n184 205.571
R4153 avdd.n306 avdd.n305 205.571
R4154 avdd.n295 avdd.n294 205.571
R4155 avdd.n284 avdd.n283 205.571
R4156 avdd.n273 avdd.n272 205.571
R4157 avdd.n322 avdd.n321 174.306
R4158 avdd.n323 avdd.n322 174.306
R4159 avdd.n345 avdd.n344 174.306
R4160 avdd.n346 avdd.n345 174.306
R4161 avdd.n369 avdd.n368 174.306
R4162 avdd.n370 avdd.n369 174.306
R4163 avdd.n393 avdd.n392 174.306
R4164 avdd.n394 avdd.n393 174.306
R4165 avdd.n328 avdd.n310 132.73
R4166 avdd.n351 avdd.n333 132.73
R4167 avdd.n375 avdd.n357 132.73
R4168 avdd.n399 avdd.n381 132.73
R4169 avdd.n329 avdd.n309 132.674
R4170 avdd.n352 avdd.n332 132.674
R4171 avdd.n376 avdd.n356 132.674
R4172 avdd.n400 avdd.n380 132.674
R4173 avdd.n86 avdd.n77 117.996
R4174 avdd.n75 avdd.n66 117.996
R4175 avdd.n64 avdd.n55 117.996
R4176 avdd.n53 avdd.n44 117.996
R4177 avdd.n42 avdd.n33 117.996
R4178 avdd.n31 avdd.n22 117.996
R4179 avdd.n20 avdd.n11 117.996
R4180 avdd.n9 avdd.n0 117.996
R4181 avdd.n174 avdd.n165 117.996
R4182 avdd.n163 avdd.n154 117.996
R4183 avdd.n152 avdd.n143 117.996
R4184 avdd.n141 avdd.n132 117.996
R4185 avdd.n130 avdd.n121 117.996
R4186 avdd.n119 avdd.n110 117.996
R4187 avdd.n108 avdd.n99 117.996
R4188 avdd.n97 avdd.n88 117.996
R4189 avdd.n262 avdd.n253 117.996
R4190 avdd.n251 avdd.n242 117.996
R4191 avdd.n240 avdd.n231 117.996
R4192 avdd.n229 avdd.n220 117.996
R4193 avdd.n218 avdd.n209 117.996
R4194 avdd.n207 avdd.n198 117.996
R4195 avdd.n196 avdd.n187 117.996
R4196 avdd.n185 avdd.n176 117.996
R4197 avdd.n306 avdd.n297 117.996
R4198 avdd.n295 avdd.n286 117.996
R4199 avdd.n284 avdd.n275 117.996
R4200 avdd.n273 avdd.n264 117.996
R4201 avdd.n325 avdd.n320 117.746
R4202 avdd.n325 avdd.n324 117.746
R4203 avdd.n348 avdd.n343 117.746
R4204 avdd.n348 avdd.n347 117.746
R4205 avdd.n372 avdd.n367 117.746
R4206 avdd.n372 avdd.n371 117.746
R4207 avdd.n396 avdd.n391 117.746
R4208 avdd.n396 avdd.n395 117.746
R4209 avdd.n321 avdd.n320 107.294
R4210 avdd.n323 avdd.n310 107.294
R4211 avdd.n324 avdd.n323 107.294
R4212 avdd.n321 avdd.n309 107.294
R4213 avdd.n344 avdd.n343 107.294
R4214 avdd.n346 avdd.n333 107.294
R4215 avdd.n347 avdd.n346 107.294
R4216 avdd.n344 avdd.n332 107.294
R4217 avdd.n368 avdd.n367 107.294
R4218 avdd.n370 avdd.n357 107.294
R4219 avdd.n371 avdd.n370 107.294
R4220 avdd.n368 avdd.n356 107.294
R4221 avdd.n392 avdd.n391 107.294
R4222 avdd.n394 avdd.n381 107.294
R4223 avdd.n395 avdd.n394 107.294
R4224 avdd.n392 avdd.n380 107.294
R4225 avdd.n80 avdd.n79 26.4291
R4226 avdd.n86 avdd.n78 26.4291
R4227 avdd.n69 avdd.n68 26.4291
R4228 avdd.n75 avdd.n67 26.4291
R4229 avdd.n58 avdd.n57 26.4291
R4230 avdd.n64 avdd.n56 26.4291
R4231 avdd.n47 avdd.n46 26.4291
R4232 avdd.n53 avdd.n45 26.4291
R4233 avdd.n36 avdd.n35 26.4291
R4234 avdd.n42 avdd.n34 26.4291
R4235 avdd.n25 avdd.n24 26.4291
R4236 avdd.n31 avdd.n23 26.4291
R4237 avdd.n14 avdd.n13 26.4291
R4238 avdd.n20 avdd.n12 26.4291
R4239 avdd.n3 avdd.n2 26.4291
R4240 avdd.n9 avdd.n1 26.4291
R4241 avdd.n168 avdd.n167 26.4291
R4242 avdd.n174 avdd.n166 26.4291
R4243 avdd.n157 avdd.n156 26.4291
R4244 avdd.n163 avdd.n155 26.4291
R4245 avdd.n146 avdd.n145 26.4291
R4246 avdd.n152 avdd.n144 26.4291
R4247 avdd.n135 avdd.n134 26.4291
R4248 avdd.n141 avdd.n133 26.4291
R4249 avdd.n124 avdd.n123 26.4291
R4250 avdd.n130 avdd.n122 26.4291
R4251 avdd.n113 avdd.n112 26.4291
R4252 avdd.n119 avdd.n111 26.4291
R4253 avdd.n102 avdd.n101 26.4291
R4254 avdd.n108 avdd.n100 26.4291
R4255 avdd.n91 avdd.n90 26.4291
R4256 avdd.n97 avdd.n89 26.4291
R4257 avdd.n256 avdd.n255 26.4291
R4258 avdd.n262 avdd.n254 26.4291
R4259 avdd.n245 avdd.n244 26.4291
R4260 avdd.n251 avdd.n243 26.4291
R4261 avdd.n234 avdd.n233 26.4291
R4262 avdd.n240 avdd.n232 26.4291
R4263 avdd.n223 avdd.n222 26.4291
R4264 avdd.n229 avdd.n221 26.4291
R4265 avdd.n212 avdd.n211 26.4291
R4266 avdd.n218 avdd.n210 26.4291
R4267 avdd.n201 avdd.n200 26.4291
R4268 avdd.n207 avdd.n199 26.4291
R4269 avdd.n190 avdd.n189 26.4291
R4270 avdd.n196 avdd.n188 26.4291
R4271 avdd.n179 avdd.n178 26.4291
R4272 avdd.n185 avdd.n177 26.4291
R4273 avdd.n300 avdd.n299 26.4291
R4274 avdd.n306 avdd.n298 26.4291
R4275 avdd.n289 avdd.n288 26.4291
R4276 avdd.n295 avdd.n287 26.4291
R4277 avdd.n278 avdd.n277 26.4291
R4278 avdd.n284 avdd.n276 26.4291
R4279 avdd.n267 avdd.n266 26.4291
R4280 avdd.n273 avdd.n265 26.4291
R4281 avdd.n320 avdd.n317 26.4291
R4282 avdd.n317 avdd.n313 26.4291
R4283 avdd.n312 avdd.n310 26.4291
R4284 avdd.n315 avdd.n312 26.4291
R4285 avdd.n324 avdd.n319 26.4291
R4286 avdd.n319 avdd.n315 26.4291
R4287 avdd.n311 avdd.n309 26.4291
R4288 avdd.n313 avdd.n311 26.4291
R4289 avdd.n343 avdd.n340 26.4291
R4290 avdd.n340 avdd.n336 26.4291
R4291 avdd.n335 avdd.n333 26.4291
R4292 avdd.n338 avdd.n335 26.4291
R4293 avdd.n347 avdd.n342 26.4291
R4294 avdd.n342 avdd.n338 26.4291
R4295 avdd.n334 avdd.n332 26.4291
R4296 avdd.n336 avdd.n334 26.4291
R4297 avdd.n367 avdd.n364 26.4291
R4298 avdd.n364 avdd.n360 26.4291
R4299 avdd.n359 avdd.n357 26.4291
R4300 avdd.n362 avdd.n359 26.4291
R4301 avdd.n371 avdd.n366 26.4291
R4302 avdd.n366 avdd.n362 26.4291
R4303 avdd.n358 avdd.n356 26.4291
R4304 avdd.n360 avdd.n358 26.4291
R4305 avdd.n391 avdd.n388 26.4291
R4306 avdd.n388 avdd.n384 26.4291
R4307 avdd.n383 avdd.n381 26.4291
R4308 avdd.n386 avdd.n383 26.4291
R4309 avdd.n395 avdd.n390 26.4291
R4310 avdd.n390 avdd.n386 26.4291
R4311 avdd.n382 avdd.n380 26.4291
R4312 avdd.n384 avdd.n382 26.4291
R4313 avdd.n81 avdd.n77 16.8187
R4314 avdd.n85 avdd.n84 16.8187
R4315 avdd.n70 avdd.n66 16.8187
R4316 avdd.n74 avdd.n73 16.8187
R4317 avdd.n59 avdd.n55 16.8187
R4318 avdd.n63 avdd.n62 16.8187
R4319 avdd.n48 avdd.n44 16.8187
R4320 avdd.n52 avdd.n51 16.8187
R4321 avdd.n37 avdd.n33 16.8187
R4322 avdd.n41 avdd.n40 16.8187
R4323 avdd.n26 avdd.n22 16.8187
R4324 avdd.n30 avdd.n29 16.8187
R4325 avdd.n15 avdd.n11 16.8187
R4326 avdd.n19 avdd.n18 16.8187
R4327 avdd.n4 avdd.n0 16.8187
R4328 avdd.n8 avdd.n7 16.8187
R4329 avdd.n169 avdd.n165 16.8187
R4330 avdd.n173 avdd.n172 16.8187
R4331 avdd.n158 avdd.n154 16.8187
R4332 avdd.n162 avdd.n161 16.8187
R4333 avdd.n147 avdd.n143 16.8187
R4334 avdd.n151 avdd.n150 16.8187
R4335 avdd.n136 avdd.n132 16.8187
R4336 avdd.n140 avdd.n139 16.8187
R4337 avdd.n125 avdd.n121 16.8187
R4338 avdd.n129 avdd.n128 16.8187
R4339 avdd.n114 avdd.n110 16.8187
R4340 avdd.n118 avdd.n117 16.8187
R4341 avdd.n103 avdd.n99 16.8187
R4342 avdd.n107 avdd.n106 16.8187
R4343 avdd.n92 avdd.n88 16.8187
R4344 avdd.n96 avdd.n95 16.8187
R4345 avdd.n257 avdd.n253 16.8187
R4346 avdd.n261 avdd.n260 16.8187
R4347 avdd.n246 avdd.n242 16.8187
R4348 avdd.n250 avdd.n249 16.8187
R4349 avdd.n235 avdd.n231 16.8187
R4350 avdd.n239 avdd.n238 16.8187
R4351 avdd.n224 avdd.n220 16.8187
R4352 avdd.n228 avdd.n227 16.8187
R4353 avdd.n213 avdd.n209 16.8187
R4354 avdd.n217 avdd.n216 16.8187
R4355 avdd.n202 avdd.n198 16.8187
R4356 avdd.n206 avdd.n205 16.8187
R4357 avdd.n191 avdd.n187 16.8187
R4358 avdd.n195 avdd.n194 16.8187
R4359 avdd.n180 avdd.n176 16.8187
R4360 avdd.n184 avdd.n183 16.8187
R4361 avdd.n301 avdd.n297 16.8187
R4362 avdd.n305 avdd.n304 16.8187
R4363 avdd.n290 avdd.n286 16.8187
R4364 avdd.n294 avdd.n293 16.8187
R4365 avdd.n279 avdd.n275 16.8187
R4366 avdd.n283 avdd.n282 16.8187
R4367 avdd.n268 avdd.n264 16.8187
R4368 avdd.n272 avdd.n271 16.8187
R4369 avdd.n326 avdd.n325 16.8187
R4370 avdd.t16 avdd.n326 16.8187
R4371 avdd.n322 avdd.n314 16.8187
R4372 avdd.t16 avdd.n314 16.8187
R4373 avdd.n328 avdd.n327 16.8187
R4374 avdd.n327 avdd.t16 16.8187
R4375 avdd.n349 avdd.n348 16.8187
R4376 avdd.t5 avdd.n349 16.8187
R4377 avdd.n345 avdd.n337 16.8187
R4378 avdd.t5 avdd.n337 16.8187
R4379 avdd.n351 avdd.n350 16.8187
R4380 avdd.n350 avdd.t5 16.8187
R4381 avdd.n373 avdd.n372 16.8187
R4382 avdd.t28 avdd.n373 16.8187
R4383 avdd.n369 avdd.n361 16.8187
R4384 avdd.t28 avdd.n361 16.8187
R4385 avdd.n375 avdd.n374 16.8187
R4386 avdd.n374 avdd.t28 16.8187
R4387 avdd.n397 avdd.n396 16.8187
R4388 avdd.t21 avdd.n397 16.8187
R4389 avdd.n393 avdd.n385 16.8187
R4390 avdd.t21 avdd.n385 16.8187
R4391 avdd.n399 avdd.n398 16.8187
R4392 avdd.n398 avdd.t21 16.8187
R4393 avdd.n82 avdd.n81 11.9049
R4394 avdd.n84 avdd.n83 11.9049
R4395 avdd.n71 avdd.n70 11.9049
R4396 avdd.n73 avdd.n72 11.9049
R4397 avdd.n60 avdd.n59 11.9049
R4398 avdd.n62 avdd.n61 11.9049
R4399 avdd.n49 avdd.n48 11.9049
R4400 avdd.n51 avdd.n50 11.9049
R4401 avdd.n38 avdd.n37 11.9049
R4402 avdd.n40 avdd.n39 11.9049
R4403 avdd.n27 avdd.n26 11.9049
R4404 avdd.n29 avdd.n28 11.9049
R4405 avdd.n16 avdd.n15 11.9049
R4406 avdd.n18 avdd.n17 11.9049
R4407 avdd.n5 avdd.n4 11.9049
R4408 avdd.n7 avdd.n6 11.9049
R4409 avdd.n170 avdd.n169 11.9049
R4410 avdd.n172 avdd.n171 11.9049
R4411 avdd.n159 avdd.n158 11.9049
R4412 avdd.n161 avdd.n160 11.9049
R4413 avdd.n148 avdd.n147 11.9049
R4414 avdd.n150 avdd.n149 11.9049
R4415 avdd.n137 avdd.n136 11.9049
R4416 avdd.n139 avdd.n138 11.9049
R4417 avdd.n126 avdd.n125 11.9049
R4418 avdd.n128 avdd.n127 11.9049
R4419 avdd.n115 avdd.n114 11.9049
R4420 avdd.n117 avdd.n116 11.9049
R4421 avdd.n104 avdd.n103 11.9049
R4422 avdd.n106 avdd.n105 11.9049
R4423 avdd.n93 avdd.n92 11.9049
R4424 avdd.n95 avdd.n94 11.9049
R4425 avdd.n258 avdd.n257 11.9049
R4426 avdd.n260 avdd.n259 11.9049
R4427 avdd.n247 avdd.n246 11.9049
R4428 avdd.n249 avdd.n248 11.9049
R4429 avdd.n236 avdd.n235 11.9049
R4430 avdd.n238 avdd.n237 11.9049
R4431 avdd.n225 avdd.n224 11.9049
R4432 avdd.n227 avdd.n226 11.9049
R4433 avdd.n214 avdd.n213 11.9049
R4434 avdd.n216 avdd.n215 11.9049
R4435 avdd.n203 avdd.n202 11.9049
R4436 avdd.n205 avdd.n204 11.9049
R4437 avdd.n192 avdd.n191 11.9049
R4438 avdd.n194 avdd.n193 11.9049
R4439 avdd.n181 avdd.n180 11.9049
R4440 avdd.n183 avdd.n182 11.9049
R4441 avdd.n302 avdd.n301 11.9049
R4442 avdd.n304 avdd.n303 11.9049
R4443 avdd.n291 avdd.n290 11.9049
R4444 avdd.n293 avdd.n292 11.9049
R4445 avdd.n280 avdd.n279 11.9049
R4446 avdd.n282 avdd.n281 11.9049
R4447 avdd.n269 avdd.n268 11.9049
R4448 avdd.n271 avdd.n270 11.9049
R4449 avdd.n407 avdd.t19 10.7165
R4450 avdd.n403 avdd.n402 6.48548
R4451 avdd.n403 avdd 4.8561
R4452 avdd.n83 avdd.t3 4.77693
R4453 avdd.t3 avdd.n82 4.77693
R4454 avdd.n72 avdd.t9 4.77693
R4455 avdd.t9 avdd.n71 4.77693
R4456 avdd.n61 avdd.t2 4.77693
R4457 avdd.t2 avdd.n60 4.77693
R4458 avdd.n50 avdd.t26 4.77693
R4459 avdd.t26 avdd.n49 4.77693
R4460 avdd.n39 avdd.t24 4.77693
R4461 avdd.t24 avdd.n38 4.77693
R4462 avdd.n28 avdd.t18 4.77693
R4463 avdd.t18 avdd.n27 4.77693
R4464 avdd.n17 avdd.t13 4.77693
R4465 avdd.t13 avdd.n16 4.77693
R4466 avdd.n6 avdd.t8 4.77693
R4467 avdd.t8 avdd.n5 4.77693
R4468 avdd.n171 avdd.t23 4.77693
R4469 avdd.t23 avdd.n170 4.77693
R4470 avdd.n160 avdd.t1 4.77693
R4471 avdd.t1 avdd.n159 4.77693
R4472 avdd.n149 avdd.t15 4.77693
R4473 avdd.t15 avdd.n148 4.77693
R4474 avdd.n138 avdd.t4 4.77693
R4475 avdd.t4 avdd.n137 4.77693
R4476 avdd.n127 avdd.t40 4.77693
R4477 avdd.t40 avdd.n126 4.77693
R4478 avdd.n116 avdd.t20 4.77693
R4479 avdd.t20 avdd.n115 4.77693
R4480 avdd.n105 avdd.t14 4.77693
R4481 avdd.t14 avdd.n104 4.77693
R4482 avdd.n94 avdd.t39 4.77693
R4483 avdd.t39 avdd.n93 4.77693
R4484 avdd.n259 avdd.t31 4.77693
R4485 avdd.t31 avdd.n258 4.77693
R4486 avdd.n248 avdd.t35 4.77693
R4487 avdd.t35 avdd.n247 4.77693
R4488 avdd.n237 avdd.t30 4.77693
R4489 avdd.t30 avdd.n236 4.77693
R4490 avdd.n226 avdd.t34 4.77693
R4491 avdd.t34 avdd.n225 4.77693
R4492 avdd.n215 avdd.t33 4.77693
R4493 avdd.t33 avdd.n214 4.77693
R4494 avdd.n204 avdd.t38 4.77693
R4495 avdd.t38 avdd.n203 4.77693
R4496 avdd.n193 avdd.t32 4.77693
R4497 avdd.t32 avdd.n192 4.77693
R4498 avdd.n182 avdd.t36 4.77693
R4499 avdd.t36 avdd.n181 4.77693
R4500 avdd.n303 avdd.t11 4.77693
R4501 avdd.t11 avdd.n302 4.77693
R4502 avdd.n292 avdd.t0 4.77693
R4503 avdd.t0 avdd.n291 4.77693
R4504 avdd.n281 avdd.t12 4.77693
R4505 avdd.t12 avdd.n280 4.77693
R4506 avdd.n270 avdd.t7 4.77693
R4507 avdd.t7 avdd.n269 4.77693
R4508 avdd.n406 avdd 3.12119
R4509 avdd.n405 avdd 3.12119
R4510 avdd.n404 avdd 3.12119
R4511 avdd avdd.n296 2.22787
R4512 avdd avdd.n274 2.22787
R4513 avdd.n10 avdd.n9 1.5505
R4514 avdd.n21 avdd.n20 1.5505
R4515 avdd.n32 avdd.n31 1.5505
R4516 avdd.n43 avdd.n42 1.5505
R4517 avdd.n54 avdd.n53 1.5505
R4518 avdd.n65 avdd.n64 1.5505
R4519 avdd.n76 avdd.n75 1.5505
R4520 avdd.n87 avdd.n86 1.5505
R4521 avdd.n98 avdd.n97 1.5505
R4522 avdd.n109 avdd.n108 1.5505
R4523 avdd.n120 avdd.n119 1.5505
R4524 avdd.n131 avdd.n130 1.5505
R4525 avdd.n142 avdd.n141 1.5505
R4526 avdd.n153 avdd.n152 1.5505
R4527 avdd.n164 avdd.n163 1.5505
R4528 avdd.n175 avdd.n174 1.5505
R4529 avdd.n186 avdd.n185 1.5505
R4530 avdd.n197 avdd.n196 1.5505
R4531 avdd.n208 avdd.n207 1.5505
R4532 avdd.n219 avdd.n218 1.5505
R4533 avdd.n230 avdd.n229 1.5505
R4534 avdd.n241 avdd.n240 1.5505
R4535 avdd.n252 avdd.n251 1.5505
R4536 avdd.n263 avdd.n262 1.5505
R4537 avdd.n274 avdd.n273 1.5505
R4538 avdd.n285 avdd.n284 1.5505
R4539 avdd.n296 avdd.n295 1.5505
R4540 avdd.n307 avdd.n306 1.5505
R4541 avdd.n354 avdd 1.38748
R4542 avdd.n378 avdd.n354 1.25871
R4543 avdd.n402 avdd.n378 1.25871
R4544 avdd.n87 avdd 1.24296
R4545 avdd.n76 avdd 1.24296
R4546 avdd.n65 avdd 1.24296
R4547 avdd.n54 avdd 1.24296
R4548 avdd.n43 avdd 1.24296
R4549 avdd.n32 avdd 1.24296
R4550 avdd.n21 avdd 1.24296
R4551 avdd.n10 avdd 1.24296
R4552 avdd.n175 avdd 1.24296
R4553 avdd.n164 avdd 1.24296
R4554 avdd.n153 avdd 1.24296
R4555 avdd.n142 avdd 1.24296
R4556 avdd.n131 avdd 1.24296
R4557 avdd.n120 avdd 1.24296
R4558 avdd.n109 avdd 1.24296
R4559 avdd.n98 avdd 1.24296
R4560 avdd.n263 avdd 1.24296
R4561 avdd.n252 avdd 1.24296
R4562 avdd.n241 avdd 1.24296
R4563 avdd.n230 avdd 1.24296
R4564 avdd.n219 avdd 1.24296
R4565 avdd.n208 avdd 1.24296
R4566 avdd.n197 avdd 1.24296
R4567 avdd.n186 avdd 1.24296
R4568 avdd.n307 avdd 1.24296
R4569 avdd.n296 avdd 1.24296
R4570 avdd.n285 avdd 1.24296
R4571 avdd.n274 avdd 1.24296
R4572 avdd avdd.n408 1.09544
R4573 avdd.n330 avdd.n329 0.645538
R4574 avdd.n353 avdd.n352 0.645538
R4575 avdd.n377 avdd.n376 0.645538
R4576 avdd.n401 avdd.n400 0.645538
R4577 avdd avdd.n87 0.492957
R4578 avdd avdd.n76 0.492957
R4579 avdd avdd.n65 0.492957
R4580 avdd avdd.n54 0.492957
R4581 avdd avdd.n43 0.492957
R4582 avdd avdd.n32 0.492957
R4583 avdd avdd.n21 0.492957
R4584 avdd avdd.n10 0.492957
R4585 avdd avdd.n175 0.492957
R4586 avdd avdd.n164 0.492957
R4587 avdd avdd.n153 0.492957
R4588 avdd avdd.n142 0.492957
R4589 avdd avdd.n131 0.492957
R4590 avdd avdd.n120 0.492957
R4591 avdd avdd.n109 0.492957
R4592 avdd avdd.n98 0.492957
R4593 avdd avdd.n263 0.492957
R4594 avdd avdd.n252 0.492957
R4595 avdd avdd.n241 0.492957
R4596 avdd avdd.n230 0.492957
R4597 avdd avdd.n219 0.492957
R4598 avdd avdd.n208 0.492957
R4599 avdd avdd.n197 0.492957
R4600 avdd avdd.n186 0.492957
R4601 avdd avdd.n307 0.492957
R4602 avdd avdd.n285 0.492957
R4603 avdd.n408 avdd.n407 0.426002
R4604 avdd.n408 avdd.n406 0.268357
R4605 avdd.n330 avdd.n308 0.265121
R4606 avdd.n353 avdd.n331 0.265121
R4607 avdd.n377 avdd.n355 0.265121
R4608 avdd.n401 avdd.n379 0.265121
R4609 avdd.n405 avdd.n404 0.148838
R4610 avdd.n404 avdd.n403 0.147954
R4611 avdd.n406 avdd.n405 0.144948
R4612 avdd.n354 avdd 0.129288
R4613 avdd.n378 avdd 0.128641
R4614 avdd.n402 avdd 0.128641
R4615 avdd.n329 avdd.n328 0.0554356
R4616 avdd.n352 avdd.n351 0.0554356
R4617 avdd.n376 avdd.n375 0.0554356
R4618 avdd.n400 avdd.n399 0.0554356
R4619 avdd avdd.n330 0.045098
R4620 avdd avdd.n353 0.045098
R4621 avdd avdd.n377 0.045098
R4622 avdd avdd.n401 0.045098
R4623 avdd.n407 avdd 0.0350686
R4624 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t11 97.2843
R4625 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t5 97.2843
R4626 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t12 24.8378
R4627 level_shifter_0.out multiplexer_0.trans_gate_m_15.ena_b 19.5921
R4628 multiplexer_0.vtrip_0.n0 multiplexer_0.trans_gate_m_8.ena 19.3217
R4629 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.n0 19.1605
R4630 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t1 18.5516
R4631 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t7 18.3731
R4632 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t4 18.1873
R4633 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t10 18.0088
R4634 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t3 16.8731
R4635 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t14 16.8731
R4636 multiplexer_0.vtrip_0.n0 multiplexer_0.vtrip_0.t16 16.8731
R4637 multiplexer_0.vtrip_0.n0 multiplexer_0.vtrip_0.t9 16.8731
R4638 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t6 16.8731
R4639 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t15 16.8731
R4640 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t8 16.5088
R4641 multiplexer_0.trans_gate_m_8.ena multiplexer_0.vtrip_0.t0 16.5088
R4642 multiplexer_0.vtrip_0.n0 multiplexer_0.vtrip_0.t2 16.5088
R4643 multiplexer_0.vtrip_0.n0 multiplexer_0.vtrip_0.t13 16.5088
R4644 multiplexer_0.trans_gate_m_15.ena_b multiplexer_0.vtrip_0.t17 16.5088
R4645 multiplexer_0.in_1011.n0 multiplexer_0.in_1011.t3 228.216
R4646 multiplexer_0.in_1011.n0 multiplexer_0.in_1011.t2 83.695
R4647 multiplexer_0.in_1011.n3 multiplexer_0.in_1011.t0 10.5295
R4648 multiplexer_0.in_1011.n3 multiplexer_0.in_1011.t1 10.5285
R4649 multiplexer_0.in_1011.n2 multiplexer_0.in_1011.n1 4.33622
R4650 multiplexer_0.in_1011.n1 multiplexer_0.in_1011.n0 1.5005
R4651 multiplexer_0.in_1011 multiplexer_0.in_1011.n3 0.872792
R4652 multiplexer_0.in_1011.n1 multiplexer_0.in_1011 0.104667
R4653 multiplexer_0.in_1011.n2 multiplexer_0.in_1011 0.0166275
R4654 multiplexer_0.in_1011 multiplexer_0.in_1011.n2 0.00984659
R4655 multiplexer_0.trans_gate_m_21.in.t5 multiplexer_0.trans_gate_m_21.in.t2 228.216
R4656 multiplexer_0.trans_gate_m_21.in.t5 multiplexer_0.trans_gate_m_21.in.t4 228.216
R4657 multiplexer_0.trans_gate_m_21.in.t5 multiplexer_0.trans_gate_m_21.in.t0 228.216
R4658 multiplexer_0.trans_gate_m_21.in.t5 multiplexer_0.trans_gate_m_21.in.t3 93.7584
R4659 multiplexer_0.trans_gate_m_21.in.t5 multiplexer_0.trans_gate_m_21.in.t1 83.695
R4660 vtrip[1].n2 vtrip[1].t2 99.4021
R4661 vtrip[1].n0 vtrip[1].t0 23.1698
R4662 vtrip[1].n1 vtrip[1].t3 17.7681
R4663 vtrip[1].n0 vtrip[1].t1 17.7475
R4664 vtrip[1].n2 vtrip[1] 5.43617
R4665 vtrip[1].n3 vtrip[1].n2 1.7055
R4666 vtrip[1].n1 vtrip[1].n0 0.572059
R4667 vtrip[1].n3 vtrip[1].n1 0.1139
R4668 vtrip[1] vtrip[1].n3 0.0378665
R4669 comp_hyst_0.net5 comp_hyst_0.net5.t2 91.2731
R4670 comp_hyst_0.net5 comp_hyst_0.net5.t0 84.6266
R4671 comp_hyst_0.net5 comp_hyst_0.net5.t1 49.1546
R4672 comp_hyst_0.net1 comp_hyst_0.net1.t3 78.9481
R4673 comp_hyst_0.net1 comp_hyst_0.net1.t2 77.4826
R4674 comp_hyst_0.net1 comp_hyst_0.net1.t1 77.4826
R4675 comp_hyst_0.net1 comp_hyst_0.net1.t0 77.4826
R4676 multiplexer_0.in_0010.n0 multiplexer_0.in_0010.t3 228.216
R4677 multiplexer_0.in_0010.n0 multiplexer_0.in_0010.t1 83.695
R4678 multiplexer_0.in_0010.n4 multiplexer_0.in_0010.t0 10.5295
R4679 multiplexer_0.in_0010.n4 multiplexer_0.in_0010.t2 10.5285
R4680 multiplexer_0.in_0010 multiplexer_0.in_0010.n3 4.90529
R4681 multiplexer_0.in_0010.n2 multiplexer_0.in_0010.n1 4.34635
R4682 multiplexer_0.in_0010.n1 multiplexer_0.in_0010.n0 1.5005
R4683 multiplexer_0.in_0010 multiplexer_0.in_0010.n4 0.872792
R4684 multiplexer_0.in_0010.n3 multiplexer_0.in_0010 0.177654
R4685 multiplexer_0.in_0010.n1 multiplexer_0.in_0010 0.104667
R4686 multiplexer_0.in_0010.n2 multiplexer_0.in_0010 0.0064902
R4687 multiplexer_0.in_0010.n3 multiplexer_0.in_0010.n2 0.00411538
R4688 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t0 227.512
R4689 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t2 99.4906
R4690 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t17 99.1756
R4691 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t1 41.0738
R4692 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t13 28.3445
R4693 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t14 22.2871
R4694 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n0 22.0358
R4695 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t10 16.8731
R4696 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t5 16.8731
R4697 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t15 16.8731
R4698 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t6 16.8731
R4699 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t3 16.8731
R4700 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t12 16.8731
R4701 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t8 16.8731
R4702 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t19 16.8731
R4703 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t16 16.5088
R4704 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t9 16.5088
R4705 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t20 16.5088
R4706 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.t11 16.5088
R4707 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t7 16.5088
R4708 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t18 16.5088
R4709 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t4 16.5088
R4710 multiplexer_0.in_0000.n0 multiplexer_0.in_0000.t1 228.216
R4711 multiplexer_0.in_0000.n0 multiplexer_0.in_0000.t2 83.695
R4712 multiplexer_0.in_0000.n3 multiplexer_0.in_0000.t0 10.5295
R4713 multiplexer_0.in_0000.n3 multiplexer_0.in_0000.t3 10.5285
R4714 multiplexer_0.in_0000 multiplexer_0.in_0000.n2 5.93817
R4715 multiplexer_0.in_0000 multiplexer_0.in_0000.n0 1.60467
R4716 multiplexer_0.in_0000 multiplexer_0.in_0000.n3 0.872792
R4717 multiplexer_0.in_0000.n2 multiplexer_0.in_0000 0.471654
R4718 multiplexer_0.in_0000.n1 multiplexer_0.in_0000 0.414042
R4719 multiplexer_0.in_0000.n1 multiplexer_0.in_0000 0.0140417
R4720 multiplexer_0.in_0000.n2 multiplexer_0.in_0000.n1 0.0101154
R4721 vin.n0 vin.t2 228.216
R4722 vin.n0 vin.t0 228.216
R4723 comp_hyst_0.vin vin.t4 101.106
R4724 vin.n0 vin.t1 83.695
R4725 vin.n0 vin.t3 83.695
R4726 vin.n0 comp_hyst_0.vin 32.334
R4727 multiplexer_0.in_1001.n0 multiplexer_0.in_1001.t2 228.216
R4728 multiplexer_0.in_1001.n0 multiplexer_0.in_1001.t1 83.695
R4729 multiplexer_0.in_1001.n2 multiplexer_0.in_1001.t0 10.5295
R4730 multiplexer_0.in_1001.n2 multiplexer_0.in_1001.t3 10.5285
R4731 multiplexer_0.in_1001 multiplexer_0.in_1001.n1 2.54596
R4732 multiplexer_0.in_1001 multiplexer_0.in_1001.n0 1.60467
R4733 multiplexer_0.in_1001 multiplexer_0.in_1001.n2 0.872792
R4734 multiplexer_0.in_1001.n1 multiplexer_0.in_1001 0.3505
R4735 multiplexer_0.in_1001.n1 multiplexer_0.in_1001 0.0775833
R4736 multiplexer_0.trans_gate_m_23.in.t2 multiplexer_0.trans_gate_m_23.in.t3 228.216
R4737 multiplexer_0.trans_gate_m_23.in.t2 multiplexer_0.trans_gate_m_23.in.t4 228.216
R4738 multiplexer_0.trans_gate_m_23.in.t2 multiplexer_0.trans_gate_m_23.in.t0 228.216
R4739 multiplexer_0.trans_gate_m_23.in.t2 multiplexer_0.trans_gate_m_23.in.t1 103.584
R4740 multiplexer_0.trans_gate_m_23.in.t2 multiplexer_0.trans_gate_m_23.in.t5 83.695
R4741 level_shifter_2.out_b multiplexer_0.vtrip_2_b.t0 227.512
R4742 multiplexer_0.trans_gate_m_32.ena multiplexer_0.vtrip_2_b.t6 99.1792
R4743 level_shifter_2.out_b multiplexer_0.vtrip_2_b.t1 41.0738
R4744 multiplexer_0.trans_gate_m_32.ena multiplexer_0.vtrip_2_b.t5 31.2886
R4745 level_shifter_2.out_b multiplexer_0.trans_gate_m_32.ena 20.4328
R4746 level_shifter_2.out_b multiplexer_0.vtrip_2_b.t2 15.633
R4747 multiplexer_0.trans_gate_m_32.ena multiplexer_0.vtrip_2_b.t3 18.5516
R4748 multiplexer_0.trans_gate_m_32.ena multiplexer_0.vtrip_2_b.t7 18.5516
R4749 multiplexer_0.trans_gate_m_32.ena multiplexer_0.vtrip_2_b.t4 18.1873
R4750 vbg.n1 vbg.t2 101.106
R4751 vbg.n0 vbg.t1 8.61346
R4752 vbg.n0 vbg.t0 8.09814
R4753 vbg.n2 vbg 4.75829
R4754 vbg vbg.n2 2.0685
R4755 vbg.n1 vbg.n0 0.303134
R4756 vbg.n2 vbg.n1 0.0129802
R4757 vbg.n2 vbg 0.00103107
R4758 multiplexer_0.in_0100.n0 multiplexer_0.in_0100.t1 228.216
R4759 multiplexer_0.in_0100.n0 multiplexer_0.in_0100.t2 83.695
R4760 multiplexer_0.in_0100.n3 multiplexer_0.in_0100.t3 10.5739
R4761 multiplexer_0.in_0100.n3 multiplexer_0.in_0100.t0 10.5739
R4762 multiplexer_0.in_0100 multiplexer_0.in_0100.n2 5.1017
R4763 multiplexer_0.in_0100 multiplexer_0.in_0100.n3 2.20538
R4764 multiplexer_0.in_0100 multiplexer_0.in_0100.n0 1.60467
R4765 multiplexer_0.in_0100.n2 multiplexer_0.in_0100 0.471654
R4766 multiplexer_0.in_0100.n1 multiplexer_0.in_0100 0.414042
R4767 multiplexer_0.in_0100.n1 multiplexer_0.in_0100 0.0140417
R4768 multiplexer_0.in_0100.n2 multiplexer_0.in_0100.n1 0.0101154
R4769 multiplexer_0.in_0101.n0 multiplexer_0.in_0101.t3 228.216
R4770 multiplexer_0.in_0101.n0 multiplexer_0.in_0101.t2 83.695
R4771 multiplexer_0.in_0101.n3 multiplexer_0.in_0101.t1 10.5739
R4772 multiplexer_0.in_0101.n3 multiplexer_0.in_0101.t0 10.5739
R4773 multiplexer_0.in_0101 multiplexer_0.in_0101.n2 4.09284
R4774 multiplexer_0.in_0101 multiplexer_0.in_0101.n3 2.20538
R4775 multiplexer_0.in_0101 multiplexer_0.in_0101.n0 1.60467
R4776 multiplexer_0.in_0101.n2 multiplexer_0.in_0101 0.471654
R4777 multiplexer_0.in_0101.n1 multiplexer_0.in_0101 0.414042
R4778 multiplexer_0.in_0101.n1 multiplexer_0.in_0101 0.0140417
R4779 multiplexer_0.in_0101.n2 multiplexer_0.in_0101.n1 0.0101154
R4780 multiplexer_0.trans_gate_m_27.in.t2 multiplexer_0.trans_gate_m_27.in.t3 228.216
R4781 multiplexer_0.trans_gate_m_27.in.t2 multiplexer_0.trans_gate_m_27.in.t4 228.216
R4782 multiplexer_0.trans_gate_m_27.in.t2 multiplexer_0.trans_gate_m_27.in.t0 228.216
R4783 multiplexer_0.trans_gate_m_27.in.t2 multiplexer_0.trans_gate_m_27.in.t1 103.584
R4784 multiplexer_0.trans_gate_m_27.in.t2 multiplexer_0.trans_gate_m_27.in.t5 83.695
R4785 multiplexer_0.trans_gate_m_28.in.t1 multiplexer_0.trans_gate_m_28.in.t2 228.216
R4786 multiplexer_0.trans_gate_m_28.in.t1 multiplexer_0.trans_gate_m_28.in.t3 228.216
R4787 multiplexer_0.trans_gate_m_28.in.t1 multiplexer_0.trans_gate_m_28.in.t0 228.216
R4788 multiplexer_0.trans_gate_m_28.in.t1 multiplexer_0.trans_gate_m_28.in.t4 93.748
R4789 ena.n9 ena.t6 99.4005
R4790 ena.n11 ena.t2 99.4005
R4791 ena.n1 ena.t7 35.2949
R4792 ena.n2 ena.t7 35.2949
R4793 ena.t3 ena.n0 34.8146
R4794 ena.n3 ena.t3 34.8146
R4795 ena.n2 ena.t1 33.8377
R4796 ena.t1 ena.n1 33.8377
R4797 ena ena.t0 25.2266
R4798 ena.n8 ena.t5 20.4065
R4799 ena.n6 ena.t5 19.344
R4800 ena.n5 ena.t4 17.6981
R4801 ena.n11 ena.n10 9.6297
R4802 ena.n10 ena 3.99824
R4803 ena.n6 ena.n5 3.48479
R4804 ena.n7 ena.n6 2.7271
R4805 ena.n4 ena.n0 1.8089
R4806 ena.n4 ena.n3 1.7055
R4807 ena.n8 ena.n7 1.7055
R4808 ena.n1 ena.n0 1.07287
R4809 ena.n3 ena.n2 1.07287
R4810 ena.n10 ena 0.46101
R4811 ena.n9 ena.n8 0.373074
R4812 ena.n5 ena.n4 0.16323
R4813 ena ena.n11 0.063
R4814 ena ena.n9 0.0309688
R4815 ena.n7 ena 0.0115247
R4816 a_n5142_n1959.t1 a_n5142_n1959.t0 41.7607
R4817 multiplexer_0.vtrip_3_b.n1 multiplexer_0.vtrip_3_b.t0 227.512
R4818 multiplexer_0.vtrip_3_b.n0 multiplexer_0.vtrip_3_b.t4 99.2037
R4819 multiplexer_0.vtrip_3_b.n1 multiplexer_0.vtrip_3_b.t1 41.0738
R4820 multiplexer_0.vtrip_3_b.n1 multiplexer_0.vtrip_3_b.n0 21.0449
R4821 multiplexer_0.vtrip_3_b.n1 multiplexer_0.vtrip_3_b.t2 16.8829
R4822 multiplexer_0.vtrip_3_b.n0 multiplexer_0.vtrip_3_b.t5 16.8731
R4823 multiplexer_0.vtrip_3_b.n0 multiplexer_0.vtrip_3_b.t3 16.5088
R4824 multiplexer_0.trans_gate_m_33.in.t2 multiplexer_0.trans_gate_m_33.in.t3 228.216
R4825 multiplexer_0.trans_gate_m_33.in.t2 multiplexer_0.trans_gate_m_33.in.t4 228.216
R4826 multiplexer_0.trans_gate_m_33.in.t2 multiplexer_0.trans_gate_m_33.in.t1 228.216
R4827 multiplexer_0.trans_gate_m_33.in.t2 multiplexer_0.trans_gate_m_33.in.t0 94.7343
R4828 multiplexer_0.in_1010.n0 multiplexer_0.in_1010.t2 228.216
R4829 multiplexer_0.in_1010.n0 multiplexer_0.in_1010.t3 83.695
R4830 multiplexer_0.in_1010.n4 multiplexer_0.in_1010.t1 10.5739
R4831 multiplexer_0.in_1010.n4 multiplexer_0.in_1010.t0 10.5739
R4832 multiplexer_0.in_1010.n2 multiplexer_0.in_1010.n1 4.34635
R4833 multiplexer_0.in_1010 multiplexer_0.in_1010.n3 3.97588
R4834 multiplexer_0.in_1010 multiplexer_0.in_1010.n4 2.20538
R4835 multiplexer_0.in_1010.n1 multiplexer_0.in_1010.n0 1.5005
R4836 multiplexer_0.in_1010.n3 multiplexer_0.in_1010 0.177654
R4837 multiplexer_0.in_1010.n1 multiplexer_0.in_1010 0.104667
R4838 multiplexer_0.in_1010.n2 multiplexer_0.in_1010 0.0064902
R4839 multiplexer_0.in_1010.n3 multiplexer_0.in_1010.n2 0.00411538
R4840 comp_hyst_0.ena_b comp_hyst_0.ena_b.t1 34.5866
R4841 comp_hyst_0.ena_b comp_hyst_0.ena_b.t1 34.5866
R4842 comp_hyst_0.ena_b comp_hyst_0.ena_b.t0 33.1294
R4843 comp_hyst_0.ena_b.t0 comp_hyst_0.ena_b 33.1294
R4844 vtrip[2].n2 vtrip[2].t3 99.4021
R4845 vtrip[2].n0 vtrip[2].t2 23.1698
R4846 vtrip[2].n1 vtrip[2].t1 17.7681
R4847 vtrip[2].n0 vtrip[2].t0 17.7475
R4848 vtrip[2].n2 vtrip[2] 5.20458
R4849 vtrip[2].n3 vtrip[2].n2 1.7055
R4850 vtrip[2].n1 vtrip[2].n0 0.572059
R4851 vtrip[2].n3 vtrip[2].n1 0.1139
R4852 vtrip[2] vtrip[2].n3 0.0378665
R4853 level_shifter_2.in_b.t1 level_shifter_2.in_b.t0 229.644
R4854 level_shifter_2.in_b.t2 level_shifter_2.in_b.t1 27.1253
R4855 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.trans_gate_m_18.in.t2 228.216
R4856 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.trans_gate_m_18.in.t4 228.216
R4857 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.trans_gate_m_18.in.t1 228.216
R4858 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.trans_gate_m_18.in.t0 103.584
R4859 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.trans_gate_m_18.in.t5 83.695
R4860 multiplexer_0.in_1110.n0 multiplexer_0.in_1110.t0 228.216
R4861 multiplexer_0.in_1110.n0 multiplexer_0.in_1110.t1 83.695
R4862 multiplexer_0.in_1110.n4 multiplexer_0.in_1110.t3 10.5739
R4863 multiplexer_0.in_1110.n4 multiplexer_0.in_1110.t2 10.5739
R4864 multiplexer_0.in_1110.n2 multiplexer_0.in_1110.n1 4.34635
R4865 multiplexer_0.in_1110 multiplexer_0.in_1110.n3 3.28049
R4866 multiplexer_0.in_1110 multiplexer_0.in_1110.n4 2.20538
R4867 multiplexer_0.in_1110.n1 multiplexer_0.in_1110.n0 1.5005
R4868 multiplexer_0.in_1110.n3 multiplexer_0.in_1110 0.177654
R4869 multiplexer_0.in_1110.n1 multiplexer_0.in_1110 0.104667
R4870 multiplexer_0.in_1110.n2 multiplexer_0.in_1110 0.0064902
R4871 multiplexer_0.in_1110.n3 multiplexer_0.in_1110.n2 0.00411538
R4872 multiplexer_0.trans_gate_m_19.in.t2 multiplexer_0.trans_gate_m_19.in.t3 228.216
R4873 multiplexer_0.trans_gate_m_19.in.t2 multiplexer_0.trans_gate_m_19.in.t5 228.216
R4874 multiplexer_0.trans_gate_m_19.in.t2 multiplexer_0.trans_gate_m_19.in.t0 228.216
R4875 multiplexer_0.trans_gate_m_19.in.t2 multiplexer_0.trans_gate_m_19.in.t4 93.7584
R4876 multiplexer_0.trans_gate_m_19.in.t2 multiplexer_0.trans_gate_m_19.in.t1 83.695
R4877 multiplexer_0.in_0011.n0 multiplexer_0.in_0011.t2 228.216
R4878 multiplexer_0.in_0011.n0 multiplexer_0.in_0011.t1 83.695
R4879 multiplexer_0.in_0011.n4 multiplexer_0.in_0011.t0 10.5295
R4880 multiplexer_0.in_0011.n4 multiplexer_0.in_0011.t3 10.5285
R4881 multiplexer_0.in_0011 multiplexer_0.in_0011.n3 4.50875
R4882 multiplexer_0.in_0011.n2 multiplexer_0.in_0011.n1 4.34635
R4883 multiplexer_0.in_0011.n1 multiplexer_0.in_0011.n0 1.5005
R4884 multiplexer_0.in_0011 multiplexer_0.in_0011.n4 0.872792
R4885 multiplexer_0.in_0011.n3 multiplexer_0.in_0011 0.177654
R4886 multiplexer_0.in_0011.n1 multiplexer_0.in_0011 0.104667
R4887 multiplexer_0.in_0011.n2 multiplexer_0.in_0011 0.0064902
R4888 multiplexer_0.in_0011.n3 multiplexer_0.in_0011.n2 0.00411538
R4889 multiplexer_0.in_0111.n0 multiplexer_0.in_0111.t2 228.216
R4890 multiplexer_0.in_0111.n0 multiplexer_0.in_0111.t1 83.695
R4891 multiplexer_0.in_0111.n4 multiplexer_0.in_0111.t0 10.5295
R4892 multiplexer_0.in_0111.n4 multiplexer_0.in_0111.t3 10.5285
R4893 multiplexer_0.in_0111.n2 multiplexer_0.in_0111.n1 4.34635
R4894 multiplexer_0.in_0111 multiplexer_0.in_0111.n3 4.17122
R4895 multiplexer_0.in_0111.n1 multiplexer_0.in_0111.n0 1.5005
R4896 multiplexer_0.in_0111 multiplexer_0.in_0111.n4 0.872792
R4897 multiplexer_0.in_0111.n3 multiplexer_0.in_0111 0.177654
R4898 multiplexer_0.in_0111.n1 multiplexer_0.in_0111 0.104667
R4899 multiplexer_0.in_0111.n2 multiplexer_0.in_0111 0.0064902
R4900 multiplexer_0.in_0111.n3 multiplexer_0.in_0111.n2 0.00411538
R4901 multiplexer_0.in_1111.n0 multiplexer_0.in_1111.t1 228.216
R4902 multiplexer_0.in_1111.n0 multiplexer_0.in_1111.t0 83.695
R4903 multiplexer_0.in_1111.n4 multiplexer_0.in_1111.t2 10.5295
R4904 multiplexer_0.in_1111.n4 multiplexer_0.in_1111.t3 10.5285
R4905 multiplexer_0.in_1111.n2 multiplexer_0.in_1111.n1 4.34635
R4906 multiplexer_0.in_1111 multiplexer_0.in_1111.n3 3.28379
R4907 multiplexer_0.in_1111.n1 multiplexer_0.in_1111.n0 1.5005
R4908 multiplexer_0.in_1111 multiplexer_0.in_1111.n4 0.872792
R4909 multiplexer_0.in_1111.n3 multiplexer_0.in_1111 0.177654
R4910 multiplexer_0.in_1111.n1 multiplexer_0.in_1111 0.104667
R4911 multiplexer_0.in_1111.n2 multiplexer_0.in_1111 0.0064902
R4912 multiplexer_0.in_1111.n3 multiplexer_0.in_1111.n2 0.00411538
R4913 multiplexer_0.trans_gate_m_25.in.t2 multiplexer_0.trans_gate_m_25.in.t3 228.216
R4914 multiplexer_0.trans_gate_m_25.in.t2 multiplexer_0.trans_gate_m_25.in.t5 228.216
R4915 multiplexer_0.trans_gate_m_25.in.t2 multiplexer_0.trans_gate_m_25.in.t0 228.216
R4916 multiplexer_0.trans_gate_m_25.in.t2 multiplexer_0.trans_gate_m_25.in.t4 93.7584
R4917 multiplexer_0.trans_gate_m_25.in.t2 multiplexer_0.trans_gate_m_25.in.t1 83.695
R4918 multiplexer_0.trans_gate_m_37.in.t1 multiplexer_0.trans_gate_m_37.in.t3 228.216
R4919 multiplexer_0.trans_gate_m_37.in.t1 multiplexer_0.trans_gate_m_37.in.t4 228.216
R4920 multiplexer_0.trans_gate_m_37.in.t1 multiplexer_0.trans_gate_m_37.in.t0 228.216
R4921 multiplexer_0.trans_gate_m_37.in.t1 multiplexer_0.trans_gate_m_37.in.t2 93.748
R4922 multiplexer_0.in_1000.n0 multiplexer_0.in_1000.t1 228.216
R4923 multiplexer_0.in_1000.n0 multiplexer_0.in_1000.t2 83.695
R4924 multiplexer_0.in_1000.n3 multiplexer_0.in_1000.t3 10.5739
R4925 multiplexer_0.in_1000.n3 multiplexer_0.in_1000.t0 10.5739
R4926 multiplexer_0.in_1000 multiplexer_0.in_1000.n2 3.76983
R4927 multiplexer_0.in_1000 multiplexer_0.in_1000.n3 2.20538
R4928 multiplexer_0.in_1000 multiplexer_0.in_1000.n0 1.60467
R4929 multiplexer_0.in_1000.n2 multiplexer_0.in_1000 0.471654
R4930 multiplexer_0.in_1000.n1 multiplexer_0.in_1000 0.414042
R4931 multiplexer_0.in_1000.n1 multiplexer_0.in_1000 0.0140417
R4932 multiplexer_0.in_1000.n2 multiplexer_0.in_1000.n1 0.0101154
R4933 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.trans_gate_m_31.in.t2 228.216
R4934 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.trans_gate_m_31.in.t4 228.216
R4935 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.trans_gate_m_31.in.t1 228.216
R4936 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.trans_gate_m_31.in.t0 103.584
R4937 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.trans_gate_m_31.in.t5 83.695
R4938 multiplexer_0.in_0001.n0 multiplexer_0.in_0001.t3 228.216
R4939 multiplexer_0.in_0001.n0 multiplexer_0.in_0001.t1 83.695
R4940 multiplexer_0.in_0001.n3 multiplexer_0.in_0001.t0 10.5295
R4941 multiplexer_0.in_0001.n3 multiplexer_0.in_0001.t2 10.5285
R4942 multiplexer_0.in_0001 multiplexer_0.in_0001.n2 4.87616
R4943 multiplexer_0.in_0001 multiplexer_0.in_0001.n0 1.60467
R4944 multiplexer_0.in_0001 multiplexer_0.in_0001.n3 0.872792
R4945 multiplexer_0.in_0001.n2 multiplexer_0.in_0001 0.471654
R4946 multiplexer_0.in_0001.n1 multiplexer_0.in_0001 0.414042
R4947 multiplexer_0.in_0001.n1 multiplexer_0.in_0001 0.0140417
R4948 multiplexer_0.in_0001.n2 multiplexer_0.in_0001.n1 0.0101154
R4949 vtrip[3].n2 vtrip[3].t3 99.4021
R4950 vtrip[3].n0 vtrip[3].t0 23.1698
R4951 vtrip[3].n1 vtrip[3].t1 17.7681
R4952 vtrip[3].n0 vtrip[3].t2 17.7475
R4953 vtrip[3].n2 vtrip[3] 4.9564
R4954 vtrip[3].n3 vtrip[3].n2 1.7055
R4955 vtrip[3].n1 vtrip[3].n0 0.572059
R4956 vtrip[3].n3 vtrip[3].n1 0.1139
R4957 vtrip[3] vtrip[3].n3 0.0378665
R4958 ibias.n0 ibias.t1 83.4559
R4959 ibias.n0 ibias.t0 42.9482
R4960 ibias.n1 ibias.n0 0.118921
R4961 ibias.n1 ibias 0.0613553
R4962 ibias ibias.n1 0.0605649
R4963 level_shifter_1.in_b.t1 level_shifter_1.in_b.t0 229.644
R4964 level_shifter_1.in_b.t2 level_shifter_1.in_b.t1 27.1253
R4965 ovout.n0 ovout.t1 92.1108
R4966 ovout.n1 ovout.t0 83.8097
R4967 ovout ovout.n1 40.1875
R4968 ovout.n0 ovout.t2 30.088
R4969 ovout.n1 ovout.n0 1.79228
C0 avss a_n12654_11271# 0.092648f
C1 m4_20244_3506# m4_19223_3506# 0.216092f
C2 m4_18268_3156# m4_18268_3506# 0.213636f
C3 avss a_n8898_4089# 0.091766f
C4 a_n8362_8625# a_n8362_7869# 0.307869f
C5 avss a_n8898_2577# 0.091766f
C6 avss a_n8898_n1203# 0.079716f
C7 avss a_n15874_309# 0.499272f
C8 a_n5142_5979# avss 0.509006f
C9 ena avdd 0.103522f
C10 multiplexer_0.in_0100 avdd 0.76049f
C11 avss multiplexer_0.in_1111 3.34253f
C12 avss a_n8898_14673# 0.094511f
C13 multiplexer_0.in_0100 multiplexer_0.vtrip_0_b 0.139372f
C14 a_n8898_1821# multiplexer_0.in_1110 0.445207f
C15 avss vtrip[2] 2.04916f
C16 avss a_n15874_13917# 0.499272f
C17 a_n8898_11649# a_n8362_11649# 0.406481f
C18 m4_18268_3506# m4_18268_4659# 0.099027f
C19 avss a_n12118_3711# 0.092648f
C20 a_n12654_10515# a_n12654_9759# 0.307869f
C21 avss a_n12654_n1203# 0.079716f
C22 dvdd comp_hyst_0.net4 30.420599f
C23 a_n5142_10515# avss 0.499272f
C24 dvdd ibias 4.8744f
C25 a_n8362_4845# multiplexer_0.in_0101 0.368184f
C26 a_n8898_13161# a_n8898_13917# 0.307869f
C27 avdd multiplexer_0.in_0011 0.6701f
C28 a_n12118_14295# a_n12654_15051# 0.307869f
C29 m4_19156_3156# m4_19223_3506# 0.249242f
C30 ovout comp_hyst_0.net4 0.385987f
C31 avss a_n12118_9759# 0.092648f
C32 a_n15874_10893# avss 0.499272f
C33 avss a_n5142_n1581# 0.499272f
C34 m4_18268_3156# m4_18268_4659# 0.012147f
C35 multiplexer_0.vtrip_0_b multiplexer_0.in_0011 0.44284f
C36 avdd multiplexer_0.in_0001 0.7344f
C37 a_n8898_10893# a_n8362_10893# 0.406481f
C38 a_n8898_4845# a_n8898_4089# 0.307869f
C39 a_n12654_3711# a_n12654_4467# 0.307869f
C40 ibias vtrip[0] 0.098883f
C41 a_n8362_7113# avss 0.092648f
C42 avss a_n5142_14295# 0.497909f
C43 a_n8898_8625# avss 0.092648f
C44 multiplexer_0.vtrip_0_b multiplexer_0.in_0001 0.144247f
C45 a_n12118_2199# avss 0.092648f
C46 avss a_n12654_8247# 0.092648f
C47 a_n15874_5601# a_n15874_4845# 0.307869f
C48 a_n5142_11271# a_n5142_12027# 0.307869f
C49 multiplexer_0.in_1111 multiplexer_0.in_1101 0.828785f
C50 a_n12654_4467# a_n12654_5223# 0.307869f
C51 a_n12654_n69# avss 0.079556f
C52 avss a_n8898_13161# 0.092648f
C53 a_n15874_8625# avss 0.499272f
C54 a_n12654_13539# a_n12654_14295# 0.307869f
C55 a_n12654_4467# a_n12118_4467# 0.406481f
C56 a_n12654_14295# a_n12118_14295# 0.406481f
C57 vtrip[1] vtrip[2] 2.74924f
C58 avss a_n12654_12783# 0.092648f
C59 multiplexer_0.in_1100 multiplexer_0.in_1001 0.02196f
C60 avdd multiplexer_0.in_1111 0.616136f
C61 avss a_n12654_9759# 0.092648f
C62 avss a_n12654_n825# 0.079566f
C63 a_n8898_7869# avss 0.092648f
C64 a_n8362_13161# a_n8362_13917# 0.307869f
C65 a_n12118_13539# a_n12654_13539# 0.406481f
C66 avdd vtrip[2] 0.206522f
C67 avss a_n8898_5601# 0.091766f
C68 multiplexer_0.in_0110 multiplexer_0.in_0000 0.01504f
C69 avss a_n12654_n1959# 0.727504f
C70 a_n12118_13539# a_n12118_14295# 0.307869f
C71 multiplexer_0.vtrip_0_b multiplexer_0.in_1111 0.463847f
C72 multiplexer_0.in_1110 multiplexer_0.in_1111 1.60188f
C73 a_n5142_n825# a_n5142_n1581# 0.307869f
C74 ovout dvdd 1.53391f
C75 ena comp_hyst_0.net5 1.53335f
C76 a_n8898_12405# a_n8898_13161# 0.307869f
C77 dvdd vtrip[0] 5.49537f
C78 a_n12654_5223# a_n12118_5223# 0.406481f
C79 a_n12118_9003# a_n12654_9003# 0.406481f
C80 a_n8898_8625# a_n8898_9381# 0.307869f
C81 multiplexer_0.in_1010 avss 2.8365f
C82 a_n12654_8247# a_n12118_8247# 0.406481f
C83 a_n12118_4467# a_n12118_5223# 0.307869f
C84 a_n8898_n69# avss 0.079556f
C85 avss a_n15874_12405# 0.499272f
C86 multiplexer_0.in_0110 avss 3.40355f
C87 a_n8898_n69# a_n8898_n447# 0.647081f
C88 a_n12654_12027# a_n12118_12027# 0.406481f
C89 a_n15874_7869# a_n15874_8625# 0.307869f
C90 avss a_n8898_n825# 0.079566f
C91 avdd a_n5142_14295# 0.374182f
C92 a_n15874_n1203# a_n15874_n1959# 0.307869f
C93 a_n12118_11271# avss 0.092648f
C94 a_n12654_687# avss 0.079556f
C95 a_n12654_11271# a_n12654_12027# 0.307869f
C96 a_n8898_n825# a_n8898_n447# 0.647081f
C97 a_n8898_n69# a_n8898_309# 0.647081f
C98 a_n8898_6357# a_n8898_5601# 0.307869f
C99 a_n12118_2199# a_n12654_1821# 0.307869f
C100 a_n12654_10515# avss 0.092648f
C101 a_n12118_7491# avss 0.092648f
C102 a_n12654_5979# avss 0.092648f
C103 a_n15874_6357# avss 0.499272f
C104 avss a_n8898_10137# 0.092648f
C105 a_n8898_4845# a_n8898_5601# 0.307869f
C106 a_n12118_10515# a_n12118_9759# 0.307869f
C107 a_n8362_12405# a_n8362_13161# 0.307869f
C108 ena comp_hyst_0.net4 0.84133f
C109 a_n8898_4089# multiplexer_0.in_1000 0.445207f
C110 a_n8362_8625# voltage_divider_0.51 0.307869f
C111 ena comp_hyst_0.net1 0.02159f
C112 multiplexer_0.in_1010 multiplexer_0.in_0111 0.930813f
C113 avss a_n8898_13917# 0.092648f
C114 avss multiplexer_0.in_0000 4.60989f
C115 ena ibias 0.657792f
C116 avss vtrip[3] 2.52607f
C117 multiplexer_0.in_0110 multiplexer_0.in_0111 1.93292f
C118 a_n5142_687# multiplexer_0.in_1111 0.368184f
C119 a_n12118_7491# a_n12118_6735# 0.307869f
C120 a_n15874_10893# a_n15874_11649# 0.307869f
C121 a_n8898_687# avss 0.079556f
C122 multiplexer_0.in_1010 avdd 0.744222f
C123 multiplexer_0.in_0100 multiplexer_0.in_0101 1.4247f
C124 a_n12118_7491# a_n12118_8247# 0.307869f
C125 multiplexer_0.in_1010 multiplexer_0.vtrip_0_b 0.490932f
C126 a_n12654_13539# a_n12654_12783# 0.307869f
C127 multiplexer_0.in_0110 avdd 0.659561f
C128 comp_hyst_0.ena_b comp_hyst_0.net5 2.09269f
C129 a_n8898_9381# a_n8898_10137# 0.307869f
C130 avss a_n12654_2955# 0.092648f
C131 multiplexer_0.in_1010 multiplexer_0.in_1110 0.01934f
C132 a_n12654_1443# avss 0.079556f
C133 avss a_n8898_n447# 0.079556f
C134 avss multiplexer_0.vtrip_1_b 10.115201f
C135 a_n8898_687# a_n8898_309# 0.647081f
C136 a_n15874_n447# a_n15874_309# 0.307869f
C137 a_n15874_4089# a_n15874_3333# 0.307869f
C138 multiplexer_0.in_0110 multiplexer_0.vtrip_0_b 0.639496f
C139 avss a_n15874_1821# 0.499272f
C140 a_n12654_n69# a_n12654_309# 0.647081f
C141 avss a_n8898_n1959# 0.727504f
C142 multiplexer_0.in_1010 multiplexer_0.in_1011 2.36311f
C143 dvdd ena 5.53155f
C144 avss a_n8898_309# 0.079556f
C145 a_n12654_12027# a_n12654_12783# 0.307869f
C146 a_n8898_3333# a_n8898_4089# 0.307869f
C147 a_n8898_3333# a_n8898_2577# 0.307869f
C148 a_n15874_10137# a_n15874_9381# 0.307869f
C149 a_n15874_6357# a_n15874_7113# 0.307869f
C150 avss a_n8898_12405# 0.092648f
C151 m4_19323_4656# m4_20044_4656# 0.248819f
C152 avss a_n12118_6735# 0.092648f
C153 ena vtrip[0] 0.314015f
C154 a_n8898_10893# a_n8898_10137# 0.307869f
C155 vtrip[3] vtrip[1] 0.374288f
C156 a_n8898_7113# a_n8362_7113# 0.406481f
C157 avdd multiplexer_0.in_0000 0.720712f
C158 a_n12118_10515# a_n12118_11271# 0.307869f
C159 a_n12654_7491# a_n12654_6735# 0.307869f
C160 a_n5142_13539# a_n5142_14295# 0.307869f
C161 a_n12654_2199# a_n12118_2199# 0.406481f
C162 a_n8898_6357# avss 0.091766f
C163 avss a_n12118_8247# 0.092648f
C164 voltage_divider_0.51 a_n8362_10137# 0.307869f
C165 a_n8898_9381# avss 0.092648f
C166 a_n12118_10515# a_n12654_10515# 0.406481f
C167 vtrip[3] avdd 0.325136f
C168 a_n8898_1443# avss 0.092791f
C169 multiplexer_0.in_0000 multiplexer_0.vtrip_0_b 0.139331f
C170 comp_hyst_0.ena_b comp_hyst_0.net4 0.014856f
C171 avss a_n5142_n825# 0.499272f
C172 avss multiplexer_0.in_0111 3.37409f
C173 comp_hyst_0.net2 comp_hyst_0.net5 0.14482f
C174 a_n15874_7869# avss 0.499272f
C175 avss multiplexer_0.in_1101 3.55535f
C176 a_n15874_12405# a_n15874_11649# 0.307869f
C177 a_n15874_4089# a_n15874_4845# 0.307869f
C178 a_n8898_4845# avss 0.092648f
C179 avss vtrip[1] 1.94321f
C180 a_n5142_5979# multiplexer_0.in_0101 0.058289f
C181 comp_hyst_0.ena_b ibias 0.812575f
C182 a_n8898_7113# a_n8898_7869# 0.307869f
C183 avss a_n5142_n69# 0.499272f
C184 multiplexer_0.vtrip_1_b vtrip[1] 0.158005f
C185 avss a_n8898_11649# 0.092648f
C186 avss a_n15874_2577# 0.499272f
C187 multiplexer_0.in_1010 multiplexer_0.in_1000 1.21062f
C188 avss avdd 1.62977p
C189 avss a_n12654_1821# 0.094199f
C190 a_n12654_687# a_n12654_309# 0.647081f
C191 a_n15874_1821# a_n15874_2577# 0.307869f
C192 a_n12654_n69# a_n12654_n447# 0.647081f
C193 avdd multiplexer_0.vtrip_1_b 10.187099f
C194 a_n15874_7113# avss 0.499272f
C195 m4_19323_4656# m4_19223_3506# 0.213636f
C196 a_n12654_1443# a_n12654_1821# 0.647081f
C197 a_n12118_9003# a_n12118_9759# 0.307869f
C198 avss multiplexer_0.vtrip_0_b 15.788701f
C199 a_n15874_309# a_n15874_1065# 0.307869f
C200 a_n8362_10893# a_n8362_10137# 0.307869f
C201 multiplexer_0.in_0110 multiplexer_0.in_1000 0.013534f
C202 avss a_n8898_10893# 0.092648f
C203 multiplexer_0.in_0100 multiplexer_0.in_0010 0.018099f
C204 a_n8898_8625# a_n8362_8625# 0.406481f
C205 avss multiplexer_0.in_1110 2.8304f
C206 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_0_b 0.705777f
C207 a_n15874_13917# a_n15874_13161# 0.307869f
C208 a_n12654_n825# a_n12654_n447# 0.647081f
C209 avss a_n12654_4467# 0.092648f
C210 a_n5142_10515# a_n5142_9759# 0.307869f
C211 a_n8898_11649# a_n8898_12405# 0.307869f
C212 dvdd vtrip[2] 3.75907f
C213 avss multiplexer_0.in_1011 3.00943f
C214 a_n12118_10515# avss 0.092648f
C215 a_n8898_687# a_n8898_1065# 0.647081f
C216 comp_hyst_0.net2 comp_hyst_0.net4 1.09495f
C217 dvdd comp_hyst_0.ena_b 2.6983f
C218 a_n8898_13161# a_n8362_13161# 0.406481f
C219 a_n8362_7113# a_n8362_7869# 0.307869f
C220 avss a_n12654_13539# 0.092648f
C221 avss a_n12118_14295# 0.092648f
C222 a_n5142_n825# a_n5142_n69# 0.307869f
C223 avss a_n8898_1065# 0.079556f
C224 vtrip[0] vtrip[2] 0.582855f
C225 multiplexer_0.in_0010 multiplexer_0.in_0011 2.38759f
C226 ovout comp_hyst_0.ena_b 0.525947f
C227 multiplexer_0.in_1100 a_n8898_2577# 0.445207f
C228 avdd multiplexer_0.in_0111 0.713663f
C229 m4_18268_3506# m4_19223_3506# 0.119924f
C230 avdd multiplexer_0.in_1101 0.704774f
C231 avss a_n15874_11649# 0.499272f
C232 avdd vtrip[1] 0.163671f
C233 multiplexer_0.in_0010 multiplexer_0.in_0001 0.856098f
C234 avss a_n12118_5223# 0.092648f
C235 multiplexer_0.vtrip_0_b multiplexer_0.in_0111 0.442759f
C236 a_n15874_7869# a_n15874_7113# 0.307869f
C237 avss a_n12654_309# 0.079556f
C238 a_n8898_7869# a_n8362_7869# 0.406481f
C239 a_n8898_3333# multiplexer_0.in_1010 0.445207f
C240 a_n8898_1443# multiplexer_0.in_1110 0.363116f
C241 multiplexer_0.vtrip_0_b multiplexer_0.in_1101 0.142054f
C242 avss a_n12654_12027# 0.092648f
C243 a_n8898_14673# a_n8362_13917# 0.307869f
C244 a_n8362_11649# a_n8362_12405# 0.307869f
C245 multiplexer_0.in_1010 multiplexer_0.in_1001 1.33401f
C246 a_n15874_10893# a_n15874_10137# 0.307869f
C247 multiplexer_0.in_1110 multiplexer_0.in_1101 1.19158f
C248 a_n8898_5601# multiplexer_0.in_0101 0.445207f
C249 avss a_n5142_12783# 0.499272f
C250 avss a_n15874_n1203# 0.499272f
C251 a_n8898_11649# a_n8898_10893# 0.307869f
C252 a_n12654_14295# a_n12654_15051# 0.307869f
C253 avdd multiplexer_0.vtrip_0_b 16.2951f
C254 m4_20044_3156# m4_20044_4656# 0.013296f
C255 avss multiplexer_0.in_1000 3.15058f
C256 multiplexer_0.in_1101 multiplexer_0.in_1011 0.313342f
C257 multiplexer_0.in_1110 avdd 0.652379f
C258 multiplexer_0.in_1010 multiplexer_0.in_0101 0.018772f
C259 a_n15874_5601# a_n15874_6357# 0.307869f
C260 a_n12654_n1581# a_n12654_n1203# 0.647081f
C261 avss a_n5142_687# 0.499272f
C262 dvdd comp_hyst_0.net2 0.550694f
C263 a_n12654_687# a_n12654_1065# 0.647081f
C264 a_n15874_13917# a_n15874_14673# 0.307869f
C265 a_n8898_1443# a_n8898_1065# 0.647081f
C266 multiplexer_0.in_1110 multiplexer_0.vtrip_0_b 0.450869f
C267 a_n8898_7113# avss 0.092648f
C268 avdd multiplexer_0.in_1011 0.836774f
C269 multiplexer_0.in_0100 multiplexer_0.in_0011 0.977996f
C270 multiplexer_0.in_0110 multiplexer_0.in_0101 1.83216f
C271 a_n12654_2199# avss 0.092648f
C272 a_n12654_2199# a_n12654_2955# 0.307869f
C273 avss a_n5142_13539# 0.499272f
C274 ovout comp_hyst_0.net2 1.14594f
C275 a_n5142_10515# a_n5142_11271# 0.307869f
C276 a_n12118_3711# a_n12118_2955# 0.307869f
C277 multiplexer_0.vtrip_0_b multiplexer_0.in_1011 0.504824f
C278 a_n8898_n1581# a_n8898_n1203# 0.647081f
C279 a_n12118_13539# a_n12118_12783# 0.307869f
C280 m4_18268_3156# m4_19156_3156# 0.186835f
C281 m4_20244_3506# m4_20044_3156# 0.122517f
C282 multiplexer_0.in_0100 multiplexer_0.in_0001 0.401107f
C283 multiplexer_0.in_1110 multiplexer_0.in_1011 0.207497f
C284 avss a_n5142_12027# 0.499272f
C285 dvdd m1_21598_448# 0.089427f
C286 a_n15874_12405# a_n15874_13161# 0.307869f
C287 avss a_n15874_n447# 0.499272f
C288 a_n8362_11649# a_n8362_10893# 0.307869f
C289 a_n12118_12027# a_n12118_12783# 0.307869f
C290 a_n8898_1821# a_n8898_2577# 0.307869f
C291 avss a_n12654_n447# 0.079556f
C292 multiplexer_0.in_1000 multiplexer_0.in_0111 1.1086f
C293 a_n15874_5601# avss 0.499272f
C294 a_n5142_5979# multiplexer_0.in_0100 0.671846f
C295 a_n8898_14673# a_n8898_15051# 0.647081f
C296 a_n12654_8247# a_n12654_9003# 0.307869f
C297 multiplexer_0.in_0000 a_n5142_9759# 0.316468f
C298 a_n8898_6357# a_n8898_7113# 0.307869f
C299 a_n8362_8625# avss 0.092648f
C300 vbg comp_hyst_0.net5 0.019445f
C301 multiplexer_0.in_0011 multiplexer_0.in_0001 0.595097f
C302 a_n8898_3333# avss 0.091766f
C303 ena vtrip[2] 0.366221f
C304 a_n12118_2199# a_n12118_2955# 0.307869f
C305 a_n12654_n1959# a_n12654_n1581# 0.647081f
C306 avss a_n12654_1065# 0.079556f
C307 avss multiplexer_0.in_1001 2.85342f
C308 avss ibias 0.011481f
C309 avdd multiplexer_0.in_1000 0.890406f
C310 avss a_n12118_9003# 0.092648f
C311 a_n5142_n69# a_n5142_687# 0.307869f
C312 a_n12654_1443# a_n12654_1065# 0.647081f
C313 avss a_n8362_13161# 0.092648f
C314 m4_19156_3156# m4_20044_3156# 0.186835f
C315 comp_hyst_0.ena_b ena 2.60102f
C316 multiplexer_0.in_1010 multiplexer_0.in_1100 0.678237f
C317 a_n12654_9759# a_n12654_9003# 0.307869f
C318 multiplexer_0.vtrip_0_b multiplexer_0.in_1000 0.140088f
C319 a_n8362_7869# avss 0.092648f
C320 a_n12654_5979# a_n12654_6735# 0.307869f
C321 a_n5142_5979# multiplexer_0.in_0011 0.313133f
C322 avss multiplexer_0.in_0101 3.35968f
C323 avss a_n5142_9759# 0.499272f
C324 a_n12654_5979# a_n12118_5979# 0.406481f
C325 a_n12654_2199# a_n12654_1821# 0.307869f
C326 dvdd vtrip[3] 2.30283f
C327 a_n12118_3711# a_n12654_3711# 0.406481f
C328 a_n8362_4845# avss 0.092648f
C329 multiplexer_0.in_1011 multiplexer_0.in_1000 0.027407f
C330 a_n8898_10137# a_n8362_10137# 0.406481f
C331 multiplexer_0.in_0100 a_n8362_7113# 0.316468f
C332 avss a_n15874_13161# 0.499272f
C333 avss a_n15874_3333# 0.499272f
C334 avss a_n15874_1065# 0.499272f
C335 vbg comp_hyst_0.net4 1.89072f
C336 vtrip[3] vtrip[0] 0.585873f
C337 a_n12118_3711# a_n12118_4467# 0.307869f
C338 a_n15874_8625# a_n15874_9381# 0.307869f
C339 a_n12118_9003# a_n12118_8247# 0.307869f
C340 vbg comp_hyst_0.net1 1.36357f
C341 avss dvdd 0.303163f
C342 a_n12654_7491# a_n12654_8247# 0.307869f
C343 multiplexer_0.in_1001 multiplexer_0.in_0111 0.31628f
C344 a_n15874_1821# a_n15874_1065# 0.307869f
C345 a_n12654_12783# a_n12118_12783# 0.406481f
C346 a_n8898_13917# a_n8362_13917# 0.406481f
C347 comp_hyst_0.net2 ena 0.032097f
C348 avss a_n15874_10137# 0.499272f
C349 avss a_n12654_6735# 0.092648f
C350 avss vtrip[0] 1.54546f
C351 avdd multiplexer_0.in_1001 0.895583f
C352 ibias avdd 0.103351f
C353 multiplexer_0.in_0111 multiplexer_0.in_0101 0.516055f
C354 a_n12118_5979# avss 0.092648f
C355 avss a_n8362_10137# 0.092648f
C356 multiplexer_0.vtrip_0_b multiplexer_0.in_1001 0.141427f
C357 multiplexer_0.in_0010 multiplexer_0.in_0000 0.748575f
C358 a_n8362_4845# a_n8898_4845# 0.406481f
C359 multiplexer_0.in_1110 multiplexer_0.in_1001 0.010731f
C360 avss multiplexer_0.in_1100 2.55289f
C361 a_n15874_4845# avss 0.499272f
C362 avss a_n8362_13917# 0.092648f
C363 avdd multiplexer_0.in_0101 0.797181f
C364 a_n5142_13539# a_n5142_12783# 0.307869f
C365 multiplexer_0.in_0110 multiplexer_0.in_0100 0.667137f
C366 multiplexer_0.in_1001 multiplexer_0.in_1011 0.660397f
C367 vbg dvdd 0.113302f
C368 avss a_n12654_n1581# 0.079868f
C369 multiplexer_0.vtrip_0_b multiplexer_0.in_0101 0.142315f
C370 a_n12654_6735# a_n12118_6735# 0.406481f
C371 a_n15874_2577# a_n15874_3333# 0.307869f
C372 dvdd vtrip[1] 3.94954f
C373 a_n5142_12027# a_n5142_12783# 0.307869f
C374 a_n12118_5979# a_n12118_6735# 0.307869f
C375 a_n5142_11271# avss 0.499272f
C376 a_n15874_n447# a_n15874_n1203# 0.307869f
C377 avss a_n15874_14673# 0.807141f
C378 multiplexer_0.in_0010 avss 4.2278f
C379 avss a_n12654_9003# 0.092648f
C380 dvdd avdd 0.213896f
C381 a_n12118_7491# a_n12654_7491# 0.406481f
C382 avss a_n12118_2955# 0.092648f
C383 vtrip[0] vtrip[1] 3.22357f
C384 a_n12654_2955# a_n12118_2955# 0.406481f
C385 multiplexer_0.in_0110 multiplexer_0.in_0011 1.4217f
C386 multiplexer_0.in_0100 multiplexer_0.in_0000 0.028175f
C387 avdd vtrip[0] 0.208605f
C388 multiplexer_0.in_1100 multiplexer_0.in_1101 1.47135f
C389 avss a_n8898_n1581# 0.079868f
C390 vtrip[3] ena 0.396701f
C391 multiplexer_0.vtrip_0_b vtrip[0] 0.158005f
C392 comp_hyst_0.ena_b comp_hyst_0.net2 0.570255f
C393 avss a_n8362_12405# 0.092648f
C394 multiplexer_0.in_1001 multiplexer_0.in_1000 1.92146f
C395 a_n12654_n825# a_n12654_n1203# 0.647081f
C396 comp_hyst_0.net5 comp_hyst_0.net4 0.078978f
C397 a_n8898_n1959# a_n8898_n1581# 0.647081f
C398 a_n12654_5979# a_n12654_5223# 0.307869f
C399 multiplexer_0.in_1100 avdd 0.655998f
C400 comp_hyst_0.net5 comp_hyst_0.net1 2.80231f
C401 avss a_n12654_15051# 0.742147f
C402 a_n12118_11271# a_n12118_12027# 0.307869f
C403 avss a_n8898_15051# 0.727504f
C404 avss a_n8898_1821# 0.091766f
C405 ibias comp_hyst_0.net5 0.720333f
C406 avss a_n15874_9381# 0.499272f
C407 a_n5142_5979# multiplexer_0.in_0110 0.309559f
C408 a_n15874_4089# avss 0.499272f
C409 avss ena 8.227719f
C410 a_n12654_9759# a_n12118_9759# 0.406481f
C411 multiplexer_0.in_0100 avss 3.71413f
C412 multiplexer_0.in_1100 multiplexer_0.vtrip_0_b 0.138847f
C413 voltage_divider_0.51 avss 0.092648f
C414 a_n12118_11271# a_n12654_11271# 0.406481f
C415 a_n8898_n825# a_n8898_n1203# 0.647081f
C416 multiplexer_0.in_1000 multiplexer_0.in_0101 0.366948f
C417 avss a_n12118_12783# 0.092648f
C418 multiplexer_0.in_1110 multiplexer_0.in_1100 0.956898f
C419 a_n12654_10515# a_n12654_11271# 0.307869f
C420 a_n12654_7491# avss 0.092648f
C421 a_n8362_4845# multiplexer_0.in_1000 0.316468f
C422 a_n8898_12405# a_n8362_12405# 0.406481f
C423 multiplexer_0.in_0000 multiplexer_0.in_0001 1.29723f
C424 m4_20244_3506# m4_20044_4656# 0.213636f
C425 a_n8898_8625# a_n8898_7869# 0.307869f
C426 multiplexer_0.in_0010 avdd 0.660581f
C427 avss a_n8362_11649# 0.092648f
C428 multiplexer_0.in_1100 multiplexer_0.in_1011 0.977944f
C429 avss a_n12654_14295# 0.092648f
C430 multiplexer_0.in_0010 multiplexer_0.vtrip_0_b 0.466038f
C431 avss a_n12654_3711# 0.092648f
C432 a_n12654_3711# a_n12654_2955# 0.307869f
C433 avss multiplexer_0.in_0011 3.46624f
C434 a_n12118_5979# a_n12118_5223# 0.307869f
C435 avss a_n8362_10893# 0.092648f
C436 avss a_n12118_13539# 0.092648f
C437 m4_19323_4656# m4_18268_4659# 0.449761f
C438 avss a_n12654_5223# 0.092648f
C439 comp_hyst_0.net1 comp_hyst_0.net4 0.063495f
C440 dvdd comp_hyst_0.net5 0.623848f
C441 a_n8898_1443# a_n8898_1821# 0.307869f
C442 a_n8898_6357# multiplexer_0.in_0100 0.445207f
C443 ibias comp_hyst_0.net4 0.049422f
C444 avss multiplexer_0.in_0001 3.89824f
C445 avss a_n12118_4467# 0.092648f
C446 a_n8898_14673# a_n8898_13917# 0.307869f
C447 a_n8898_9381# voltage_divider_0.51 0.406481f
C448 avss a_n12118_12027# 0.092648f
C449 avss a_n15874_n1959# 0.807141f
C450 ovout comp_hyst_0.net5 0.038309f
C451 vtrip[3] vtrip[2] 2.12757f
C452 ena vtrip[1] 0.370864f
C453 vbg dvss 11.814878f
C454 ovout dvss 4.14261f
C455 ibias dvss 9.874781f
C456 ena dvss 20.711246f
C457 vtrip[3] dvss 7.803799f
C458 vtrip[2] dvss 9.231338f
C459 vtrip[1] dvss 9.753779f
C460 vtrip[0] dvss 10.507146f
C461 avss dvss 0.406581p
C462 dvdd dvss 1.216993p
C463 avdd dvss 2.03821p
C464 m4_20044_3156# dvss 0.49052f $ **FLOATING
C465 m4_19156_3156# dvss 0.34028f $ **FLOATING
C466 m4_18268_3156# dvss 0.496944f $ **FLOATING
C467 m4_20244_3506# dvss 0.332279f $ **FLOATING
C468 m4_19223_3506# dvss 0.2996f $ **FLOATING
C469 m4_18268_3506# dvss 0.388269f $ **FLOATING
C470 m4_20044_4656# dvss 0.610775f $ **FLOATING
C471 m4_19323_4656# dvss 0.296713f $ **FLOATING
C472 m4_18268_4659# dvss 0.695734f $ **FLOATING
C473 m1_21598_448# dvss 4.41071f $ **FLOATING
C474 comp_hyst_0.net1 dvss 7.30358f
C475 comp_hyst_0.net5 dvss 29.79036f
C476 comp_hyst_0.net2 dvss 7.539189f
C477 comp_hyst_0.ena_b dvss 16.282839f
C478 comp_hyst_0.net4 dvss 12.0192f
C479 multiplexer_0.vtrip_1_b dvss 24.398848f
C480 multiplexer_0.vtrip_0_b dvss 26.01862f
C481 a_n8898_n1959# dvss 0.503897f
C482 a_n12654_n1959# dvss 0.503897f
C483 a_n8898_n1581# dvss 0.503897f
C484 a_n12654_n1581# dvss 0.503897f
C485 a_n15874_n1959# dvss 0.506846f
C486 a_n5142_n1581# dvss 0.506846f
C487 a_n8898_n1203# dvss 0.503897f
C488 a_n12654_n1203# dvss 0.503897f
C489 a_n8898_n825# dvss 0.503897f
C490 a_n12654_n825# dvss 0.503897f
C491 a_n15874_n1203# dvss 0.506846f
C492 a_n5142_n825# dvss 0.506846f
C493 a_n8898_n447# dvss 0.503897f
C494 a_n12654_n447# dvss 0.503897f
C495 a_n8898_n69# dvss 0.503897f
C496 a_n12654_n69# dvss 0.503897f
C497 a_n15874_n447# dvss 0.506846f
C498 a_n5142_n69# dvss 0.506846f
C499 a_n8898_309# dvss 0.503897f
C500 a_n12654_309# dvss 0.503897f
C501 a_n8898_687# dvss 0.503897f
C502 a_n12654_687# dvss 0.503897f
C503 a_n15874_309# dvss 0.506846f
C504 a_n5142_687# dvss 0.506846f
C505 a_n8898_1065# dvss 0.503897f
C506 a_n12654_1065# dvss 0.503897f
C507 a_n8898_1443# dvss 0.506785f
C508 a_n12654_1443# dvss 0.503897f
C509 a_n15874_1065# dvss 0.506846f
C510 multiplexer_0.in_1111 dvss 1.823567f
C511 a_n12654_1821# dvss 0.507092f
C512 multiplexer_0.in_1110 dvss 2.124716f
C513 a_n8898_1821# dvss 0.506846f
C514 a_n15874_1821# dvss 0.506846f
C515 multiplexer_0.in_1101 dvss 1.810742f
C516 a_n12118_2199# dvss 0.506846f
C517 a_n12654_2199# dvss 0.506846f
C518 multiplexer_0.in_1100 dvss 1.583226f
C519 a_n8898_2577# dvss 0.506846f
C520 a_n15874_2577# dvss 0.506846f
C521 multiplexer_0.in_1011 dvss 2.71753f
C522 a_n12118_2955# dvss 0.506846f
C523 a_n12654_2955# dvss 0.506846f
C524 multiplexer_0.in_1010 dvss 2.890666f
C525 a_n8898_3333# dvss 0.506846f
C526 a_n15874_3333# dvss 0.506846f
C527 multiplexer_0.in_1001 dvss 1.689299f
C528 a_n12118_3711# dvss 0.506846f
C529 a_n12654_3711# dvss 0.506846f
C530 multiplexer_0.in_1000 dvss 2.181204f
C531 a_n8898_4089# dvss 0.506846f
C532 a_n15874_4089# dvss 0.506846f
C533 multiplexer_0.in_0111 dvss 1.826988f
C534 a_n12118_4467# dvss 0.506846f
C535 a_n12654_4467# dvss 0.506846f
C536 a_n8362_4845# dvss 0.506846f
C537 a_n8898_4845# dvss 0.506846f
C538 a_n15874_4845# dvss 0.506846f
C539 multiplexer_0.in_0110 dvss 1.901118f
C540 a_n12118_5223# dvss 0.506846f
C541 a_n12654_5223# dvss 0.506846f
C542 multiplexer_0.in_0101 dvss 2.265734f
C543 a_n8898_5601# dvss 0.506846f
C544 a_n15874_5601# dvss 0.506846f
C545 a_n5142_5979# dvss 0.508215f
C546 a_n12118_5979# dvss 0.506846f
C547 a_n12654_5979# dvss 0.506846f
C548 multiplexer_0.in_0100 dvss 2.550706f
C549 a_n8898_6357# dvss 0.506846f
C550 a_n15874_6357# dvss 0.506846f
C551 multiplexer_0.in_0011 dvss 2.577745f
C552 a_n12118_6735# dvss 0.506846f
C553 a_n12654_6735# dvss 0.506846f
C554 a_n8362_7113# dvss 0.506846f
C555 a_n8898_7113# dvss 0.506846f
C556 a_n15874_7113# dvss 0.506846f
C557 multiplexer_0.in_0010 dvss 3.263069f
C558 a_n12118_7491# dvss 0.506846f
C559 a_n12654_7491# dvss 0.506846f
C560 a_n8362_7869# dvss 0.506846f
C561 a_n8898_7869# dvss 0.506846f
C562 a_n15874_7869# dvss 0.506846f
C563 multiplexer_0.in_0001 dvss 1.934929f
C564 a_n12118_8247# dvss 0.506846f
C565 a_n12654_8247# dvss 0.506846f
C566 a_n8362_8625# dvss 0.506846f
C567 a_n8898_8625# dvss 0.506846f
C568 a_n15874_8625# dvss 0.506846f
C569 multiplexer_0.in_0000 dvss 2.276361f
C570 a_n12118_9003# dvss 0.506846f
C571 a_n12654_9003# dvss 0.506846f
C572 voltage_divider_0.51 dvss 0.506846f
C573 a_n8898_9381# dvss 0.506846f
C574 a_n15874_9381# dvss 0.506846f
C575 a_n5142_9759# dvss 0.506846f
C576 a_n12118_9759# dvss 0.506846f
C577 a_n12654_9759# dvss 0.506846f
C578 a_n8362_10137# dvss 0.506846f
C579 a_n8898_10137# dvss 0.506846f
C580 a_n15874_10137# dvss 0.506846f
C581 a_n5142_10515# dvss 0.506846f
C582 a_n12118_10515# dvss 0.506846f
C583 a_n12654_10515# dvss 0.506846f
C584 a_n8362_10893# dvss 0.506846f
C585 a_n8898_10893# dvss 0.506846f
C586 a_n15874_10893# dvss 0.506846f
C587 a_n5142_11271# dvss 0.506846f
C588 a_n12118_11271# dvss 0.506846f
C589 a_n12654_11271# dvss 0.506846f
C590 a_n8362_11649# dvss 0.506846f
C591 a_n8898_11649# dvss 0.506846f
C592 a_n15874_11649# dvss 0.506846f
C593 a_n5142_12027# dvss 0.506846f
C594 a_n12118_12027# dvss 0.506846f
C595 a_n12654_12027# dvss 0.506846f
C596 a_n8362_12405# dvss 0.506846f
C597 a_n8898_12405# dvss 0.506846f
C598 a_n15874_12405# dvss 0.506846f
C599 a_n5142_12783# dvss 0.506846f
C600 a_n12118_12783# dvss 0.506846f
C601 a_n12654_12783# dvss 0.506846f
C602 a_n8362_13161# dvss 0.506846f
C603 a_n8898_13161# dvss 0.506846f
C604 a_n15874_13161# dvss 0.506846f
C605 a_n5142_13539# dvss 0.506846f
C606 a_n12118_13539# dvss 0.506846f
C607 a_n12654_13539# dvss 0.506846f
C608 a_n8362_13917# dvss 0.506846f
C609 a_n8898_13917# dvss 0.506846f
C610 a_n15874_13917# dvss 0.506846f
C611 a_n5142_14295# dvss 0.506846f
C612 a_n8898_14673# dvss 0.507092f
C613 a_n12118_14295# dvss 0.506846f
C614 a_n12654_14295# dvss 0.506846f
C615 a_n8898_15051# dvss 0.503897f
C616 a_n12654_15051# dvss 0.507092f
C617 a_n15874_14673# dvss 0.506846f
C618 level_shifter_1.in_b.t0 dvss 0.045956f
C619 level_shifter_1.in_b.t1 dvss 2.92589f
C620 level_shifter_1.in_b.t2 dvss 1.52816f
C621 ibias.t1 dvss 0.020303f
C622 ibias.t0 dvss 0.151424f
C623 ibias.n0 dvss 0.560183f
C624 ibias.n1 dvss 0.010762f
C625 vtrip[3].t0 dvss 0.971899f
C626 vtrip[3].t2 dvss 0.646085f
C627 vtrip[3].n0 dvss 1.65578f
C628 vtrip[3].t1 dvss 0.61254f
C629 vtrip[3].n1 dvss 2.1534f
C630 vtrip[3].t3 dvss 0.041792f
C631 vtrip[3].n2 dvss 0.765388f
C632 vtrip[3].n3 dvss 0.344f
C633 multiplexer_0.in_0001.t3 dvss 0.020428f
C634 multiplexer_0.in_0001.t1 dvss 0.019952f
C635 multiplexer_0.in_0001.n0 dvss 0.174642f
C636 multiplexer_0.in_0001.n1 dvss 0.04807f
C637 multiplexer_0.in_0001.n2 dvss 0.368274f
C638 multiplexer_0.in_0001.t2 dvss 0.078554f
C639 multiplexer_0.in_0001.t0 dvss 0.078563f
C640 multiplexer_0.in_0001.n3 dvss 1.76738f
C641 multiplexer_0.trans_gate_m_31.in.t3 dvss 3.27656f
C642 multiplexer_0.trans_gate_m_31.in.t2 dvss 0.024921f
C643 multiplexer_0.trans_gate_m_31.in.t0 dvss 0.02434f
C644 multiplexer_0.trans_gate_m_31.in.t4 dvss 0.024921f
C645 multiplexer_0.trans_gate_m_31.in.t5 dvss 0.02434f
C646 multiplexer_0.trans_gate_m_31.in.t1 dvss 0.024921f
C647 multiplexer_0.in_1000.t1 dvss 0.011299f
C648 multiplexer_0.in_1000.t2 dvss 0.011036f
C649 multiplexer_0.in_1000.n0 dvss 0.096602f
C650 multiplexer_0.in_1000.n1 dvss 0.02659f
C651 multiplexer_0.in_1000.n2 dvss 0.145999f
C652 multiplexer_0.in_1000.t3 dvss 0.043538f
C653 multiplexer_0.in_1000.t0 dvss 0.043538f
C654 multiplexer_0.in_1000.n3 dvss 1.48678f
C655 multiplexer_0.trans_gate_m_37.in.t1 dvss 3.05134f
C656 multiplexer_0.trans_gate_m_37.in.t0 dvss 0.037383f
C657 multiplexer_0.trans_gate_m_37.in.t3 dvss 0.037383f
C658 multiplexer_0.trans_gate_m_37.in.t4 dvss 0.037383f
C659 multiplexer_0.trans_gate_m_37.in.t2 dvss 0.036512f
C660 multiplexer_0.trans_gate_m_25.in.t2 dvss 2.73241f
C661 multiplexer_0.trans_gate_m_25.in.t5 dvss 0.033834f
C662 multiplexer_0.trans_gate_m_25.in.t4 dvss 0.033046f
C663 multiplexer_0.trans_gate_m_25.in.t3 dvss 0.033834f
C664 multiplexer_0.trans_gate_m_25.in.t1 dvss 0.033046f
C665 multiplexer_0.trans_gate_m_25.in.t0 dvss 0.033834f
C666 multiplexer_0.in_1111.t1 dvss 0.01764f
C667 multiplexer_0.in_1111.t0 dvss 0.017229f
C668 multiplexer_0.in_1111.n0 dvss 0.148902f
C669 multiplexer_0.in_1111.n1 dvss 0.093583f
C670 multiplexer_0.in_1111.n2 dvss 0.333201f
C671 multiplexer_0.in_1111.n3 dvss 0.228318f
C672 multiplexer_0.in_1111.t3 dvss 0.067836f
C673 multiplexer_0.in_1111.t2 dvss 0.067844f
C674 multiplexer_0.in_1111.n4 dvss 1.52623f
C675 multiplexer_0.in_0111.t2 dvss 0.015206f
C676 multiplexer_0.in_0111.t1 dvss 0.014851f
C677 multiplexer_0.in_0111.n0 dvss 0.12835f
C678 multiplexer_0.in_0111.n1 dvss 0.080666f
C679 multiplexer_0.in_0111.n2 dvss 0.287213f
C680 multiplexer_0.in_0111.n3 dvss 0.315379f
C681 multiplexer_0.in_0111.t3 dvss 0.058473f
C682 multiplexer_0.in_0111.t0 dvss 0.05848f
C683 multiplexer_0.in_0111.n4 dvss 1.31558f
C684 multiplexer_0.in_0011.t2 dvss 0.025975f
C685 multiplexer_0.in_0011.t1 dvss 0.025369f
C686 multiplexer_0.in_0011.n0 dvss 0.21925f
C687 multiplexer_0.in_0011.n1 dvss 0.137796f
C688 multiplexer_0.in_0011.n2 dvss 0.490621f
C689 multiplexer_0.in_0011.n3 dvss 0.675355f
C690 multiplexer_0.in_0011.t3 dvss 0.099885f
C691 multiplexer_0.in_0011.t0 dvss 0.099896f
C692 multiplexer_0.in_0011.n4 dvss 2.24729f
C693 multiplexer_0.trans_gate_m_19.in.t2 dvss 2.82663f
C694 multiplexer_0.trans_gate_m_19.in.t5 dvss 0.035001f
C695 multiplexer_0.trans_gate_m_19.in.t4 dvss 0.034185f
C696 multiplexer_0.trans_gate_m_19.in.t3 dvss 0.035001f
C697 multiplexer_0.trans_gate_m_19.in.t1 dvss 0.034185f
C698 multiplexer_0.trans_gate_m_19.in.t0 dvss 0.035001f
C699 multiplexer_0.in_1110.n0 dvss 0.083691f
C700 multiplexer_0.in_1110.n1 dvss 0.052599f
C701 multiplexer_0.in_1110.n2 dvss 0.187277f
C702 multiplexer_0.in_1110.n3 dvss 0.122179f
C703 multiplexer_0.in_1110.t3 dvss 0.038204f
C704 multiplexer_0.in_1110.t2 dvss 0.038204f
C705 multiplexer_0.in_1110.n4 dvss 1.30461f
C706 multiplexer_0.trans_gate_m_18.in.t3 dvss 3.27656f
C707 multiplexer_0.trans_gate_m_18.in.t2 dvss 0.024921f
C708 multiplexer_0.trans_gate_m_18.in.t0 dvss 0.02434f
C709 multiplexer_0.trans_gate_m_18.in.t4 dvss 0.024921f
C710 multiplexer_0.trans_gate_m_18.in.t5 dvss 0.02434f
C711 multiplexer_0.trans_gate_m_18.in.t1 dvss 0.024921f
C712 level_shifter_2.in_b.t0 dvss 0.045956f
C713 level_shifter_2.in_b.t1 dvss 2.92589f
C714 level_shifter_2.in_b.t2 dvss 1.52816f
C715 vtrip[2].t2 dvss 1.21331f
C716 vtrip[2].t0 dvss 0.806564f
C717 vtrip[2].n0 dvss 2.06705f
C718 vtrip[2].t1 dvss 0.764687f
C719 vtrip[2].n1 dvss 2.68828f
C720 vtrip[2].t3 dvss 0.052172f
C721 vtrip[2].n2 dvss 1.29487f
C722 vtrip[2].n3 dvss 0.429445f
C723 comp_hyst_0.ena_b.t1 dvss 0.363228f
C724 comp_hyst_0.ena_b.t0 dvss 0.340927f
C725 multiplexer_0.in_1010.t2 dvss 0.016668f
C726 multiplexer_0.in_1010.t3 dvss 0.01628f
C727 multiplexer_0.in_1010.n0 dvss 0.140696f
C728 multiplexer_0.in_1010.n1 dvss 0.088425f
C729 multiplexer_0.in_1010.n2 dvss 0.314839f
C730 multiplexer_0.in_1010.n3 dvss 0.298874f
C731 multiplexer_0.in_1010.t1 dvss 0.064225f
C732 multiplexer_0.in_1010.t0 dvss 0.064225f
C733 multiplexer_0.in_1010.n4 dvss 2.19323f
C734 multiplexer_0.trans_gate_m_33.in.t2 dvss 4.15315f
C735 multiplexer_0.trans_gate_m_33.in.t4 dvss 0.036927f
C736 multiplexer_0.trans_gate_m_33.in.t3 dvss 0.036927f
C737 multiplexer_0.trans_gate_m_33.in.t0 dvss 0.036067f
C738 multiplexer_0.trans_gate_m_33.in.t1 dvss 0.036927f
C739 multiplexer_0.vtrip_3_b.n0 dvss 5.71966f
C740 multiplexer_0.vtrip_3_b.n1 dvss 3.47039f
C741 multiplexer_0.vtrip_3_b.t4 dvss 0.061793f
C742 multiplexer_0.vtrip_3_b.t3 dvss 0.798611f
C743 multiplexer_0.vtrip_3_b.t5 dvss 0.829687f
C744 multiplexer_0.vtrip_3_b.t1 dvss 0.091521f
C745 multiplexer_0.vtrip_3_b.t0 dvss 0.048044f
C746 multiplexer_0.vtrip_3_b.t2 dvss 0.880296f
C747 a_n5142_n1959.t0 dvss 0.900602f
C748 a_n5142_n1959.t1 dvss 2.3994f
C749 ena.t5 dvss 0.484358f
C750 ena.n0 dvss 0.269051f
C751 ena.t3 dvss 0.304155f
C752 ena.t7 dvss 0.310806f
C753 ena.n1 dvss 0.422771f
C754 ena.t1 dvss 0.293114f
C755 ena.n2 dvss 0.422771f
C756 ena.n3 dvss 0.265961f
C757 ena.n4 dvss 0.253884f
C758 ena.t4 dvss 0.313176f
C759 ena.n5 dvss 1.0283f
C760 ena.n6 dvss 0.459201f
C761 ena.n7 dvss 0.120055f
C762 ena.n8 dvss 0.355583f
C763 ena.t6 dvss 0.021453f
C764 ena.n9 dvss 0.061353f
C765 ena.n10 dvss 5.0478f
C766 ena.t2 dvss 0.021334f
C767 ena.n11 dvss 2.97276f
C768 ena.t0 dvss 0.535271f
C769 multiplexer_0.trans_gate_m_28.in.t1 dvss 2.76528f
C770 multiplexer_0.trans_gate_m_28.in.t0 dvss 0.033878f
C771 multiplexer_0.trans_gate_m_28.in.t2 dvss 0.033878f
C772 multiplexer_0.trans_gate_m_28.in.t4 dvss 0.033089f
C773 multiplexer_0.trans_gate_m_28.in.t3 dvss 0.033878f
C774 multiplexer_0.trans_gate_m_27.in.t2 dvss 3.18019f
C775 multiplexer_0.trans_gate_m_27.in.t3 dvss 0.024188f
C776 multiplexer_0.trans_gate_m_27.in.t1 dvss 0.023624f
C777 multiplexer_0.trans_gate_m_27.in.t4 dvss 0.024188f
C778 multiplexer_0.trans_gate_m_27.in.t5 dvss 0.023624f
C779 multiplexer_0.trans_gate_m_27.in.t0 dvss 0.024188f
C780 multiplexer_0.in_0101.t3 dvss 0.012096f
C781 multiplexer_0.in_0101.t2 dvss 0.011814f
C782 multiplexer_0.in_0101.n0 dvss 0.103412f
C783 multiplexer_0.in_0101.n1 dvss 0.028464f
C784 multiplexer_0.in_0101.n2 dvss 0.166739f
C785 multiplexer_0.in_0101.t1 dvss 0.046607f
C786 multiplexer_0.in_0101.t0 dvss 0.046607f
C787 multiplexer_0.in_0101.n3 dvss 1.5916f
C788 multiplexer_0.in_0100.t1 dvss 0.012875f
C789 multiplexer_0.in_0100.t2 dvss 0.012575f
C790 multiplexer_0.in_0100.n0 dvss 0.110071f
C791 multiplexer_0.in_0100.n1 dvss 0.030297f
C792 multiplexer_0.in_0100.n2 dvss 0.242516f
C793 multiplexer_0.in_0100.t3 dvss 0.049609f
C794 multiplexer_0.in_0100.t0 dvss 0.049609f
C795 multiplexer_0.in_0100.n3 dvss 1.6941f
C796 vbg.t1 dvss 0.574937f
C797 vbg.t0 dvss 0.536153f
C798 vbg.n0 dvss 1.25899f
C799 vbg.t2 dvss 0.011064f
C800 vbg.n1 dvss 0.154849f
C801 vbg.n2 dvss 0.150024f
C802 multiplexer_0.trans_gate_m_32.ena dvss 10.5835f
C803 level_shifter_2.out_b dvss 3.3275f
C804 multiplexer_0.vtrip_2_b.t1 dvss 0.081691f
C805 multiplexer_0.vtrip_2_b.t0 dvss 0.042884f
C806 multiplexer_0.vtrip_2_b.t5 dvss 0.776964f
C807 multiplexer_0.vtrip_2_b.t7 dvss 0.806147f
C808 multiplexer_0.vtrip_2_b.t6 dvss 0.055259f
C809 multiplexer_0.vtrip_2_b.t4 dvss 0.776962f
C810 multiplexer_0.vtrip_2_b.t3 dvss 0.806147f
C811 multiplexer_0.vtrip_2_b.t2 dvss 0.742982f
C812 multiplexer_0.trans_gate_m_23.in.t2 dvss 3.27656f
C813 multiplexer_0.trans_gate_m_23.in.t3 dvss 0.024921f
C814 multiplexer_0.trans_gate_m_23.in.t1 dvss 0.02434f
C815 multiplexer_0.trans_gate_m_23.in.t4 dvss 0.024921f
C816 multiplexer_0.trans_gate_m_23.in.t5 dvss 0.02434f
C817 multiplexer_0.trans_gate_m_23.in.t0 dvss 0.024921f
C818 multiplexer_0.in_1001.t2 dvss 0.015872f
C819 multiplexer_0.in_1001.t1 dvss 0.015502f
C820 multiplexer_0.in_1001.n0 dvss 0.135692f
C821 multiplexer_0.in_1001.n1 dvss 0.13812f
C822 multiplexer_0.in_1001.t3 dvss 0.061035f
C823 multiplexer_0.in_1001.t0 dvss 0.061041f
C824 multiplexer_0.in_1001.n2 dvss 1.3732f
C825 vin.n0 dvss 2.10253f
C826 comp_hyst_0.vin dvss 5.03028f
C827 vin.t2 dvss 0.012759f
C828 vin.t1 dvss 0.012462f
C829 vin.t4 dvss 0.016742f
C830 vin.t0 dvss 0.012759f
C831 vin.t3 dvss 0.012462f
C832 multiplexer_0.in_0000.t1 dvss 0.023325f
C833 multiplexer_0.in_0000.t2 dvss 0.022782f
C834 multiplexer_0.in_0000.n0 dvss 0.199413f
C835 multiplexer_0.in_0000.n1 dvss 0.054889f
C836 multiplexer_0.in_0000.n2 dvss 0.547631f
C837 multiplexer_0.in_0000.t3 dvss 0.089697f
C838 multiplexer_0.in_0000.t0 dvss 0.089707f
C839 multiplexer_0.in_0000.n3 dvss 2.01807f
C840 multiplexer_0.vtrip_0_b.n0 dvss 10.2891f
C841 multiplexer_0.vtrip_0_b.t1 dvss 0.08376f
C842 multiplexer_0.vtrip_0_b.t0 dvss 0.04397f
C843 multiplexer_0.vtrip_0_b.t17 dvss 0.056646f
C844 multiplexer_0.vtrip_0_b.t9 dvss 0.73089f
C845 multiplexer_0.vtrip_0_b.t5 dvss 0.759332f
C846 multiplexer_0.vtrip_0_b.t16 dvss 0.73089f
C847 multiplexer_0.vtrip_0_b.t10 dvss 0.759332f
C848 multiplexer_0.vtrip_0_b.t2 dvss 0.057901f
C849 multiplexer_0.vtrip_0_b.t4 dvss 0.73089f
C850 multiplexer_0.vtrip_0_b.t19 dvss 0.759332f
C851 multiplexer_0.vtrip_0_b.t13 dvss 0.73089f
C852 multiplexer_0.vtrip_0_b.t8 dvss 0.759332f
C853 multiplexer_0.vtrip_0_b.t18 dvss 0.73089f
C854 multiplexer_0.vtrip_0_b.t12 dvss 0.759332f
C855 multiplexer_0.vtrip_0_b.t7 dvss 0.73089f
C856 multiplexer_0.vtrip_0_b.t3 dvss 0.759332f
C857 multiplexer_0.vtrip_0_b.t11 dvss 0.73089f
C858 multiplexer_0.vtrip_0_b.t6 dvss 0.759332f
C859 multiplexer_0.vtrip_0_b.t20 dvss 0.73089f
C860 multiplexer_0.vtrip_0_b.t15 dvss 0.759332f
C861 multiplexer_0.vtrip_0_b.t14 dvss 0.761802f
C862 multiplexer_0.in_0010.t3 dvss 0.028311f
C863 multiplexer_0.in_0010.t1 dvss 0.027652f
C864 multiplexer_0.in_0010.n0 dvss 0.238974f
C865 multiplexer_0.in_0010.n1 dvss 0.150192f
C866 multiplexer_0.in_0010.n2 dvss 0.534759f
C867 multiplexer_0.in_0010.n3 dvss 0.877195f
C868 multiplexer_0.in_0010.t2 dvss 0.108871f
C869 multiplexer_0.in_0010.t0 dvss 0.108883f
C870 multiplexer_0.in_0010.n4 dvss 2.44947f
C871 comp_hyst_0.net1.t3 dvss 0.046148f
C872 comp_hyst_0.net1.t0 dvss 0.04377f
C873 comp_hyst_0.net1.t1 dvss 0.04377f
C874 comp_hyst_0.net1.t2 dvss 0.04377f
C875 comp_hyst_0.net5.t2 dvss 0.0131f
C876 comp_hyst_0.net5.t1 dvss 0.068132f
C877 vtrip[1].t0 dvss 1.03496f
C878 vtrip[1].t1 dvss 0.688005f
C879 vtrip[1].n0 dvss 1.76321f
C880 vtrip[1].t3 dvss 0.652284f
C881 vtrip[1].n1 dvss 2.29313f
C882 vtrip[1].t2 dvss 0.044504f
C883 vtrip[1].n2 dvss 1.48872f
C884 vtrip[1].n3 dvss 0.36632f
C885 multiplexer_0.trans_gate_m_21.in.t5 dvss 2.82663f
C886 multiplexer_0.trans_gate_m_21.in.t4 dvss 0.035001f
C887 multiplexer_0.trans_gate_m_21.in.t3 dvss 0.034185f
C888 multiplexer_0.trans_gate_m_21.in.t2 dvss 0.035001f
C889 multiplexer_0.trans_gate_m_21.in.t1 dvss 0.034185f
C890 multiplexer_0.trans_gate_m_21.in.t0 dvss 0.035001f
C891 multiplexer_0.in_1011.t3 dvss 0.025514f
C892 multiplexer_0.in_1011.t2 dvss 0.02492f
C893 multiplexer_0.in_1011.n0 dvss 0.215366f
C894 multiplexer_0.in_1011.n1 dvss 0.134241f
C895 multiplexer_0.in_1011.n2 dvss 0.486091f
C896 multiplexer_0.in_1011.t1 dvss 0.098115f
C897 multiplexer_0.in_1011.t0 dvss 0.098127f
C898 multiplexer_0.in_1011.n3 dvss 2.20748f
C899 multiplexer_0.vtrip_0.n0 dvss 6.1358f
C900 multiplexer_0.trans_gate_m_15.ena_b dvss 11.6685f
C901 multiplexer_0.trans_gate_m_8.ena dvss 9.55242f
C902 multiplexer_0.vtrip_0.t1 dvss 1.0194f
C903 multiplexer_0.vtrip_0.t7 dvss 1.01084f
C904 multiplexer_0.vtrip_0.t11 dvss 0.066195f
C905 multiplexer_0.vtrip_0.t12 dvss 0.901404f
C906 multiplexer_0.vtrip_0.t15 dvss 0.936482f
C907 multiplexer_0.vtrip_0.t17 dvss 0.901404f
C908 multiplexer_0.vtrip_0.t6 dvss 0.936482f
C909 multiplexer_0.vtrip_0.t4 dvss 0.982498f
C910 multiplexer_0.vtrip_0.t10 dvss 0.974118f
C911 multiplexer_0.vtrip_0.t5 dvss 0.066195f
C912 multiplexer_0.vtrip_0.t0 dvss 0.901404f
C913 multiplexer_0.vtrip_0.t14 dvss 0.936482f
C914 multiplexer_0.vtrip_0.t8 dvss 0.901404f
C915 multiplexer_0.vtrip_0.t3 dvss 0.936482f
C916 multiplexer_0.vtrip_0.t13 dvss 0.901404f
C917 multiplexer_0.vtrip_0.t9 dvss 0.936482f
C918 multiplexer_0.vtrip_0.t2 dvss 0.901404f
C919 multiplexer_0.vtrip_0.t16 dvss 0.936482f
C920 level_shifter_0.out dvss 6.99673f
C921 avdd.n0 dvss 0.800453f
C922 avdd.n1 dvss 5.39489f
C923 avdd.n2 dvss 0.488536f
C924 avdd.n3 dvss 5.39489f
C925 avdd.n4 dvss 0.811075f
C926 avdd.t8 dvss 7.22231f
C927 avdd.n7 dvss 0.811075f
C928 avdd.n8 dvss 0.446622f
C929 avdd.n9 dvss 2.06399f
C930 avdd.n10 dvss 1.72384f
C931 avdd.n11 dvss 0.800453f
C932 avdd.n12 dvss 5.39489f
C933 avdd.n13 dvss 0.488536f
C934 avdd.n14 dvss 5.39489f
C935 avdd.n15 dvss 0.811075f
C936 avdd.t13 dvss 7.22231f
C937 avdd.n18 dvss 0.811075f
C938 avdd.n19 dvss 0.446622f
C939 avdd.n20 dvss 2.06399f
C940 avdd.n21 dvss 1.72384f
C941 avdd.n22 dvss 0.800453f
C942 avdd.n23 dvss 5.39489f
C943 avdd.n24 dvss 0.488536f
C944 avdd.n25 dvss 5.39489f
C945 avdd.n26 dvss 0.811075f
C946 avdd.t18 dvss 7.22231f
C947 avdd.n29 dvss 0.811075f
C948 avdd.n30 dvss 0.446622f
C949 avdd.n31 dvss 2.06399f
C950 avdd.n32 dvss 1.72384f
C951 avdd.n33 dvss 0.800453f
C952 avdd.n34 dvss 5.39489f
C953 avdd.n35 dvss 0.488536f
C954 avdd.n36 dvss 5.39489f
C955 avdd.n37 dvss 0.811075f
C956 avdd.t24 dvss 7.22231f
C957 avdd.n40 dvss 0.811075f
C958 avdd.n41 dvss 0.446622f
C959 avdd.n42 dvss 2.06399f
C960 avdd.n43 dvss 1.72384f
C961 avdd.n44 dvss 0.800453f
C962 avdd.n45 dvss 5.39489f
C963 avdd.n46 dvss 0.488536f
C964 avdd.n47 dvss 5.39489f
C965 avdd.n48 dvss 0.811075f
C966 avdd.t26 dvss 7.22231f
C967 avdd.n51 dvss 0.811075f
C968 avdd.n52 dvss 0.446622f
C969 avdd.n53 dvss 2.06399f
C970 avdd.n54 dvss 1.72384f
C971 avdd.n55 dvss 0.800453f
C972 avdd.n56 dvss 5.39489f
C973 avdd.n57 dvss 0.488536f
C974 avdd.n58 dvss 5.39489f
C975 avdd.n59 dvss 0.811075f
C976 avdd.t2 dvss 7.22231f
C977 avdd.n62 dvss 0.811075f
C978 avdd.n63 dvss 0.446622f
C979 avdd.n64 dvss 2.06399f
C980 avdd.n65 dvss 1.72384f
C981 avdd.n66 dvss 0.800453f
C982 avdd.n67 dvss 5.39489f
C983 avdd.n68 dvss 0.488536f
C984 avdd.n69 dvss 5.39489f
C985 avdd.n70 dvss 0.811075f
C986 avdd.t9 dvss 7.22231f
C987 avdd.n73 dvss 0.811075f
C988 avdd.n74 dvss 0.446622f
C989 avdd.n75 dvss 2.06399f
C990 avdd.n76 dvss 1.72384f
C991 avdd.n77 dvss 0.800453f
C992 avdd.n78 dvss 5.39489f
C993 avdd.n79 dvss 0.488536f
C994 avdd.n80 dvss 5.39489f
C995 avdd.n81 dvss 0.811075f
C996 avdd.t3 dvss 7.22231f
C997 avdd.n84 dvss 0.811075f
C998 avdd.n85 dvss 0.446622f
C999 avdd.n86 dvss 2.06399f
C1000 avdd.n87 dvss 1.72384f
C1001 avdd.n88 dvss 0.800453f
C1002 avdd.n89 dvss 5.39489f
C1003 avdd.n90 dvss 0.488536f
C1004 avdd.n91 dvss 5.39489f
C1005 avdd.n92 dvss 0.811075f
C1006 avdd.t39 dvss 7.22231f
C1007 avdd.n95 dvss 0.811075f
C1008 avdd.n96 dvss 0.446622f
C1009 avdd.n97 dvss 2.06399f
C1010 avdd.n98 dvss 1.72384f
C1011 avdd.n99 dvss 0.800453f
C1012 avdd.n100 dvss 5.39489f
C1013 avdd.n101 dvss 0.488536f
C1014 avdd.n102 dvss 5.39489f
C1015 avdd.n103 dvss 0.811075f
C1016 avdd.t14 dvss 7.22231f
C1017 avdd.n106 dvss 0.811075f
C1018 avdd.n107 dvss 0.446622f
C1019 avdd.n108 dvss 2.06399f
C1020 avdd.n109 dvss 1.72384f
C1021 avdd.n110 dvss 0.800453f
C1022 avdd.n111 dvss 5.39489f
C1023 avdd.n112 dvss 0.488536f
C1024 avdd.n113 dvss 5.39489f
C1025 avdd.n114 dvss 0.811075f
C1026 avdd.t20 dvss 7.22231f
C1027 avdd.n117 dvss 0.811075f
C1028 avdd.n118 dvss 0.446622f
C1029 avdd.n119 dvss 2.06399f
C1030 avdd.n120 dvss 1.72384f
C1031 avdd.n121 dvss 0.800453f
C1032 avdd.n122 dvss 5.39489f
C1033 avdd.n123 dvss 0.488536f
C1034 avdd.n124 dvss 5.39489f
C1035 avdd.n125 dvss 0.811075f
C1036 avdd.t40 dvss 7.22231f
C1037 avdd.n128 dvss 0.811075f
C1038 avdd.n129 dvss 0.446622f
C1039 avdd.n130 dvss 2.06399f
C1040 avdd.n131 dvss 1.72384f
C1041 avdd.n132 dvss 0.800453f
C1042 avdd.n133 dvss 5.39489f
C1043 avdd.n134 dvss 0.488536f
C1044 avdd.n135 dvss 5.39489f
C1045 avdd.n136 dvss 0.811075f
C1046 avdd.t4 dvss 7.22231f
C1047 avdd.n139 dvss 0.811075f
C1048 avdd.n140 dvss 0.446622f
C1049 avdd.n141 dvss 2.06399f
C1050 avdd.n142 dvss 1.72384f
C1051 avdd.n143 dvss 0.800453f
C1052 avdd.n144 dvss 5.39489f
C1053 avdd.n145 dvss 0.488536f
C1054 avdd.n146 dvss 5.39489f
C1055 avdd.n147 dvss 0.811075f
C1056 avdd.t15 dvss 7.22231f
C1057 avdd.n150 dvss 0.811075f
C1058 avdd.n151 dvss 0.446622f
C1059 avdd.n152 dvss 2.06399f
C1060 avdd.n153 dvss 1.72384f
C1061 avdd.n154 dvss 0.800453f
C1062 avdd.n155 dvss 5.39489f
C1063 avdd.n156 dvss 0.488536f
C1064 avdd.n157 dvss 5.39489f
C1065 avdd.n158 dvss 0.811075f
C1066 avdd.t1 dvss 7.22231f
C1067 avdd.n161 dvss 0.811075f
C1068 avdd.n162 dvss 0.446622f
C1069 avdd.n163 dvss 2.06399f
C1070 avdd.n164 dvss 1.72384f
C1071 avdd.n165 dvss 0.800453f
C1072 avdd.n166 dvss 5.39489f
C1073 avdd.n167 dvss 0.488536f
C1074 avdd.n168 dvss 5.39489f
C1075 avdd.n169 dvss 0.811075f
C1076 avdd.t23 dvss 7.22231f
C1077 avdd.n172 dvss 0.811075f
C1078 avdd.n173 dvss 0.446622f
C1079 avdd.n174 dvss 2.06399f
C1080 avdd.n175 dvss 1.72384f
C1081 avdd.n176 dvss 0.800453f
C1082 avdd.n177 dvss 5.39489f
C1083 avdd.n178 dvss 0.488536f
C1084 avdd.n179 dvss 5.39489f
C1085 avdd.n180 dvss 0.811075f
C1086 avdd.t36 dvss 7.22231f
C1087 avdd.n183 dvss 0.811075f
C1088 avdd.n184 dvss 0.446622f
C1089 avdd.n185 dvss 2.06399f
C1090 avdd.n186 dvss 1.72384f
C1091 avdd.n187 dvss 0.800453f
C1092 avdd.n188 dvss 5.39489f
C1093 avdd.n189 dvss 0.488536f
C1094 avdd.n190 dvss 5.39489f
C1095 avdd.n191 dvss 0.811075f
C1096 avdd.t32 dvss 7.22231f
C1097 avdd.n194 dvss 0.811075f
C1098 avdd.n195 dvss 0.446622f
C1099 avdd.n196 dvss 2.06399f
C1100 avdd.n197 dvss 1.72384f
C1101 avdd.n198 dvss 0.800453f
C1102 avdd.n199 dvss 5.39489f
C1103 avdd.n200 dvss 0.488536f
C1104 avdd.n201 dvss 5.39489f
C1105 avdd.n202 dvss 0.811075f
C1106 avdd.t38 dvss 7.22231f
C1107 avdd.n205 dvss 0.811075f
C1108 avdd.n206 dvss 0.446622f
C1109 avdd.n207 dvss 2.06399f
C1110 avdd.n208 dvss 1.72384f
C1111 avdd.n209 dvss 0.800453f
C1112 avdd.n210 dvss 5.39489f
C1113 avdd.n211 dvss 0.488536f
C1114 avdd.n212 dvss 5.39489f
C1115 avdd.n213 dvss 0.811075f
C1116 avdd.t33 dvss 7.22231f
C1117 avdd.n216 dvss 0.811075f
C1118 avdd.n217 dvss 0.446622f
C1119 avdd.n218 dvss 2.06399f
C1120 avdd.n219 dvss 1.72384f
C1121 avdd.n220 dvss 0.800453f
C1122 avdd.n221 dvss 5.39489f
C1123 avdd.n222 dvss 0.488536f
C1124 avdd.n223 dvss 5.39489f
C1125 avdd.n224 dvss 0.811075f
C1126 avdd.t34 dvss 7.22231f
C1127 avdd.n227 dvss 0.811075f
C1128 avdd.n228 dvss 0.446622f
C1129 avdd.n229 dvss 2.06399f
C1130 avdd.n230 dvss 1.72384f
C1131 avdd.n231 dvss 0.800453f
C1132 avdd.n232 dvss 5.39489f
C1133 avdd.n233 dvss 0.488536f
C1134 avdd.n234 dvss 5.39489f
C1135 avdd.n235 dvss 0.811075f
C1136 avdd.t30 dvss 7.22231f
C1137 avdd.n238 dvss 0.811075f
C1138 avdd.n239 dvss 0.446622f
C1139 avdd.n240 dvss 2.06399f
C1140 avdd.n241 dvss 1.72384f
C1141 avdd.n242 dvss 0.800453f
C1142 avdd.n243 dvss 5.39489f
C1143 avdd.n244 dvss 0.488536f
C1144 avdd.n245 dvss 5.39489f
C1145 avdd.n246 dvss 0.811075f
C1146 avdd.t35 dvss 7.22231f
C1147 avdd.n249 dvss 0.811075f
C1148 avdd.n250 dvss 0.446622f
C1149 avdd.n251 dvss 2.06399f
C1150 avdd.n252 dvss 1.72384f
C1151 avdd.n253 dvss 0.800453f
C1152 avdd.n254 dvss 5.39489f
C1153 avdd.n255 dvss 0.488536f
C1154 avdd.n256 dvss 5.39489f
C1155 avdd.n257 dvss 0.811075f
C1156 avdd.t31 dvss 7.22231f
C1157 avdd.n260 dvss 0.811075f
C1158 avdd.n261 dvss 0.446622f
C1159 avdd.n262 dvss 2.06399f
C1160 avdd.n263 dvss 1.72384f
C1161 avdd.n264 dvss 0.800453f
C1162 avdd.n265 dvss 5.39489f
C1163 avdd.n266 dvss 0.488536f
C1164 avdd.n267 dvss 5.39489f
C1165 avdd.n268 dvss 0.811075f
C1166 avdd.t7 dvss 7.22231f
C1167 avdd.n271 dvss 0.811075f
C1168 avdd.n272 dvss 0.446622f
C1169 avdd.n273 dvss 2.06399f
C1170 avdd.n274 dvss 3.44767f
C1171 avdd.n275 dvss 0.800453f
C1172 avdd.n276 dvss 5.39489f
C1173 avdd.n277 dvss 0.488536f
C1174 avdd.n278 dvss 5.39489f
C1175 avdd.n279 dvss 0.811075f
C1176 avdd.t12 dvss 7.22231f
C1177 avdd.n282 dvss 0.811075f
C1178 avdd.n283 dvss 0.446622f
C1179 avdd.n284 dvss 2.06399f
C1180 avdd.n285 dvss 1.72384f
C1181 avdd.n286 dvss 0.800453f
C1182 avdd.n287 dvss 5.39489f
C1183 avdd.n288 dvss 0.488536f
C1184 avdd.n289 dvss 5.39489f
C1185 avdd.n290 dvss 0.811075f
C1186 avdd.t0 dvss 7.22231f
C1187 avdd.n293 dvss 0.811075f
C1188 avdd.n294 dvss 0.446622f
C1189 avdd.n295 dvss 2.06399f
C1190 avdd.n296 dvss 3.44767f
C1191 avdd.n297 dvss 0.800453f
C1192 avdd.n298 dvss 5.39489f
C1193 avdd.n299 dvss 0.488536f
C1194 avdd.n300 dvss 5.39489f
C1195 avdd.n301 dvss 0.811075f
C1196 avdd.t11 dvss 7.22231f
C1197 avdd.n304 dvss 0.811075f
C1198 avdd.n305 dvss 0.446622f
C1199 avdd.n306 dvss 2.06399f
C1200 avdd.n307 dvss 1.72384f
C1201 avdd.t27 dvss 0.200137f
C1202 avdd.t17 dvss 0.197247f
C1203 avdd.n308 dvss 2.802f
C1204 avdd.n309 dvss 0.400052f
C1205 avdd.n310 dvss 0.400849f
C1206 avdd.n311 dvss 0.559704f
C1207 avdd.n312 dvss 0.559704f
C1208 avdd.n313 dvss 8.426219f
C1209 avdd.n314 dvss 0.495737f
C1210 avdd.n315 dvss 8.426219f
C1211 avdd.n316 dvss 0.571222f
C1212 avdd.n317 dvss 0.559704f
C1213 avdd.n318 dvss 0.571222f
C1214 avdd.n319 dvss 0.559704f
C1215 avdd.n320 dvss 0.417714f
C1216 avdd.n321 dvss 0.334854f
C1217 avdd.n322 dvss 0.290604f
C1218 avdd.n323 dvss 0.334854f
C1219 avdd.n324 dvss 0.417714f
C1220 avdd.n325 dvss 9.74957f
C1221 avdd.n326 dvss 0.811075f
C1222 avdd.t16 dvss 11.948999f
C1223 avdd.n327 dvss 0.811075f
C1224 avdd.n328 dvss 1.93421f
C1225 avdd.n329 dvss 2.93397f
C1226 avdd.n330 dvss 2.80158f
C1227 avdd.t6 dvss 0.200137f
C1228 avdd.t10 dvss 0.197247f
C1229 avdd.n331 dvss 2.802f
C1230 avdd.n332 dvss 0.400052f
C1231 avdd.n333 dvss 0.400849f
C1232 avdd.n334 dvss 0.559704f
C1233 avdd.n335 dvss 0.559704f
C1234 avdd.n336 dvss 8.426219f
C1235 avdd.n337 dvss 0.495737f
C1236 avdd.n338 dvss 8.426219f
C1237 avdd.n339 dvss 0.571222f
C1238 avdd.n340 dvss 0.559704f
C1239 avdd.n341 dvss 0.571222f
C1240 avdd.n342 dvss 0.559704f
C1241 avdd.n343 dvss 0.417714f
C1242 avdd.n344 dvss 0.334854f
C1243 avdd.n345 dvss 0.290604f
C1244 avdd.n346 dvss 0.334854f
C1245 avdd.n347 dvss 0.417714f
C1246 avdd.n348 dvss 9.74957f
C1247 avdd.n349 dvss 0.811075f
C1248 avdd.t5 dvss 11.948999f
C1249 avdd.n350 dvss 0.811075f
C1250 avdd.n351 dvss 1.93421f
C1251 avdd.n352 dvss 2.93397f
C1252 avdd.n353 dvss 2.80158f
C1253 avdd.n354 dvss 8.42617f
C1254 avdd.t37 dvss 0.200137f
C1255 avdd.t29 dvss 0.197247f
C1256 avdd.n355 dvss 2.802f
C1257 avdd.n356 dvss 0.400052f
C1258 avdd.n357 dvss 0.400849f
C1259 avdd.n358 dvss 0.559704f
C1260 avdd.n359 dvss 0.559704f
C1261 avdd.n360 dvss 8.426219f
C1262 avdd.n361 dvss 0.495737f
C1263 avdd.n362 dvss 8.426219f
C1264 avdd.n363 dvss 0.571222f
C1265 avdd.n364 dvss 0.559704f
C1266 avdd.n365 dvss 0.571222f
C1267 avdd.n366 dvss 0.559704f
C1268 avdd.n367 dvss 0.417714f
C1269 avdd.n368 dvss 0.334854f
C1270 avdd.n369 dvss 0.290604f
C1271 avdd.n370 dvss 0.334854f
C1272 avdd.n371 dvss 0.417714f
C1273 avdd.n372 dvss 9.74957f
C1274 avdd.n373 dvss 0.811075f
C1275 avdd.t28 dvss 11.948999f
C1276 avdd.n374 dvss 0.811075f
C1277 avdd.n375 dvss 1.93421f
C1278 avdd.n376 dvss 2.93397f
C1279 avdd.n377 dvss 2.80158f
C1280 avdd.n378 dvss 8.02315f
C1281 avdd.t25 dvss 0.200137f
C1282 avdd.t22 dvss 0.197247f
C1283 avdd.n379 dvss 2.802f
C1284 avdd.n380 dvss 0.400052f
C1285 avdd.n381 dvss 0.400849f
C1286 avdd.n382 dvss 0.559704f
C1287 avdd.n383 dvss 0.559704f
C1288 avdd.n384 dvss 8.426219f
C1289 avdd.n385 dvss 0.495737f
C1290 avdd.n386 dvss 8.426219f
C1291 avdd.n387 dvss 0.571222f
C1292 avdd.n388 dvss 0.559704f
C1293 avdd.n389 dvss 0.571222f
C1294 avdd.n390 dvss 0.559704f
C1295 avdd.n391 dvss 0.417714f
C1296 avdd.n392 dvss 0.334854f
C1297 avdd.n393 dvss 0.290604f
C1298 avdd.n394 dvss 0.334854f
C1299 avdd.n395 dvss 0.417714f
C1300 avdd.n396 dvss 9.74957f
C1301 avdd.n397 dvss 0.811075f
C1302 avdd.t21 dvss 11.948999f
C1303 avdd.n398 dvss 0.811075f
C1304 avdd.n399 dvss 1.93421f
C1305 avdd.n400 dvss 2.93397f
C1306 avdd.n401 dvss 2.80158f
C1307 avdd.n402 dvss 24.6949f
C1308 avdd.n403 dvss 0.105131p
C1309 avdd.n404 dvss 46.7712f
C1310 avdd.n405 dvss 46.327503f
C1311 avdd.n406 dvss 63.9731f
C1312 avdd.t19 dvss 0.873456f
C1313 avdd.n407 dvss 13.3624f
C1314 avdd.n408 dvss 0.20923p
C1315 multiplexer_0.trans_gate_m_37.out.t3 dvss 4.02134f
C1316 multiplexer_0.trans_gate_m_37.out.t5 dvss 0.036068f
C1317 multiplexer_0.trans_gate_m_37.out.t4 dvss 0.035228f
C1318 multiplexer_0.trans_gate_m_37.out.t2 dvss 0.036068f
C1319 multiplexer_0.trans_gate_m_37.out.t0 dvss 0.035228f
C1320 multiplexer_0.trans_gate_m_37.out.t1 dvss 0.036068f
C1321 multiplexer_0.trans_gate_m_32.in.t0 dvss 2.86063f
C1322 multiplexer_0.trans_gate_m_32.in.t1 dvss 0.035046f
C1323 multiplexer_0.trans_gate_m_32.in.t2 dvss 0.035046f
C1324 multiplexer_0.trans_gate_m_32.in.t4 dvss 0.035046f
C1325 multiplexer_0.trans_gate_m_32.in.t3 dvss 0.03423f
C1326 level_shifter_0.in_b.t0 dvss 0.022467f
C1327 level_shifter_0.in_b.t1 dvss 1.43043f
C1328 level_shifter_0.in_b.t2 dvss 0.7471f
C1329 vtrip[0].t1 dvss 0.855519f
C1330 vtrip[0].t0 dvss 0.568719f
C1331 vtrip[0].n0 dvss 1.45751f
C1332 vtrip[0].t3 dvss 0.539191f
C1333 vtrip[0].n1 dvss 1.89554f
C1334 vtrip[0].t2 dvss 0.036787f
C1335 vtrip[0].n2 dvss 1.6207f
C1336 vtrip[0].n3 dvss 0.302807f
C1337 multiplexer_0.in_1101.t0 dvss 0.02041f
C1338 multiplexer_0.in_1101.t1 dvss 0.019934f
C1339 multiplexer_0.in_1101.n0 dvss 0.174486f
C1340 multiplexer_0.in_1101.n1 dvss 0.048028f
C1341 multiplexer_0.in_1101.n2 dvss 0.291486f
C1342 multiplexer_0.in_1101.t3 dvss 0.078484f
C1343 multiplexer_0.in_1101.t2 dvss 0.078493f
C1344 multiplexer_0.in_1101.n3 dvss 1.7658f
C1345 multiplexer_0.in_1100.t1 dvss 0.010459f
C1346 multiplexer_0.in_1100.t2 dvss 0.010216f
C1347 multiplexer_0.in_1100.n0 dvss 0.089419f
C1348 multiplexer_0.in_1100.n1 dvss 0.024613f
C1349 multiplexer_0.in_1100.n2 dvss 0.059537f
C1350 multiplexer_0.in_1100.t3 dvss 0.040301f
C1351 multiplexer_0.in_1100.t0 dvss 0.040301f
C1352 multiplexer_0.in_1100.n3 dvss 1.37623f
C1353 multiplexer_0.vtrip_2.n0 dvss 2.12286f
C1354 multiplexer_0.trans_gate_m_20.ena_b dvss 11.0057f
C1355 level_shifter_2.out dvss 4.9667f
C1356 multiplexer_0.vtrip_2.t0 dvss 0.060235f
C1357 multiplexer_0.vtrip_2.t5 dvss 1.09443f
C1358 multiplexer_0.vtrip_2.t3 dvss 1.1353f
C1359 multiplexer_0.vtrip_2.t4 dvss 1.00389f
C1360 multiplexer_0.vtrip_2.t2 dvss 1.04296f
C1361 multiplexer_0.vtrip_2.t1 dvss 0.073735f
C1362 multiplexer_0.vtrip_2.t6 dvss 1.09421f
C1363 multiplexer_0.in_0110.t2 dvss 0.01481f
C1364 multiplexer_0.in_0110.t1 dvss 0.014465f
C1365 multiplexer_0.in_0110.n0 dvss 0.125009f
C1366 multiplexer_0.in_0110.n1 dvss 0.078566f
C1367 multiplexer_0.in_0110.n2 dvss 0.279735f
C1368 multiplexer_0.in_0110.n3 dvss 0.375647f
C1369 multiplexer_0.in_0110.t3 dvss 0.056951f
C1370 multiplexer_0.in_0110.t0 dvss 0.056957f
C1371 multiplexer_0.in_0110.n4 dvss 1.28133f
C1372 multiplexer_0.trans_gate_m_33.ena_b dvss 6.98391f
C1373 multiplexer_0.vtrip_3.n0 dvss 4.13561f
C1374 multiplexer_0.vtrip_3.t5 dvss 1.00938f
C1375 multiplexer_0.vtrip_3.t4 dvss 0.065556f
C1376 multiplexer_0.vtrip_3.t3 dvss 0.97284f
C1377 multiplexer_0.vtrip_3.t0 dvss 0.10611f
C1378 multiplexer_0.vtrip_3.t1 dvss 0.053554f
C1379 multiplexer_0.vtrip_3.t2 dvss 0.97304f
C1380 level_shifter_3.in_b.t1 dvss 0.046977f
C1381 level_shifter_3.in_b.t0 dvss 2.99091f
C1382 level_shifter_3.in_b.t2 dvss 1.56212f
C1383 comp_hyst_0.net3.t0 dvss 63.2878f
C1384 comp_hyst_0.net3.t3 dvss 0.093209f
C1385 comp_hyst_0.net3.t1 dvss 0.04075f
C1386 comp_hyst_0.net3.t2 dvss 0.078278f
C1387 dvdd.n0 dvss 0.02099f
C1388 dvdd.n1 dvss 0.123013f
C1389 dvdd.t96 dvss 0.218923f
C1390 dvdd.n3 dvss 0.140612f
C1391 dvdd.n4 dvss 0.016706f
C1392 dvdd.n5 dvss 0.017574f
C1393 dvdd.n7 dvss 0.140612f
C1394 dvdd.n8 dvss 0.017574f
C1395 dvdd.n9 dvss 0.073445f
C1396 dvdd.n10 dvss 0.109985f
C1397 dvdd.n11 dvss 0.136347f
C1398 dvdd.n12 dvss 0.02099f
C1399 dvdd.n13 dvss 0.123013f
C1400 dvdd.t109 dvss 0.218923f
C1401 dvdd.n15 dvss 0.140612f
C1402 dvdd.n16 dvss 0.016706f
C1403 dvdd.n17 dvss 0.017574f
C1404 dvdd.n19 dvss 0.140612f
C1405 dvdd.n20 dvss 0.017574f
C1406 dvdd.n21 dvss 0.073445f
C1407 dvdd.n22 dvss 0.109985f
C1408 dvdd.n23 dvss 0.136347f
C1409 dvdd.n24 dvss 0.02099f
C1410 dvdd.n25 dvss 0.123013f
C1411 dvdd.t111 dvss 0.218923f
C1412 dvdd.n27 dvss 0.140612f
C1413 dvdd.n28 dvss 0.016706f
C1414 dvdd.n29 dvss 0.017574f
C1415 dvdd.n31 dvss 0.140612f
C1416 dvdd.n32 dvss 0.017574f
C1417 dvdd.n33 dvss 0.073445f
C1418 dvdd.n34 dvss 0.109985f
C1419 dvdd.n35 dvss 0.136347f
C1420 dvdd.n36 dvss 0.02099f
C1421 dvdd.n37 dvss 0.123013f
C1422 dvdd.t92 dvss 0.218923f
C1423 dvdd.n39 dvss 0.140612f
C1424 dvdd.n40 dvss 0.016706f
C1425 dvdd.n41 dvss 0.017574f
C1426 dvdd.n43 dvss 0.140612f
C1427 dvdd.n44 dvss 0.017574f
C1428 dvdd.n45 dvss 0.073445f
C1429 dvdd.n46 dvss 0.109985f
C1430 dvdd.n47 dvss 0.136347f
C1431 dvdd.n48 dvss 0.081677f
C1432 dvdd.n49 dvss 0.623931f
C1433 dvdd.n50 dvss 2.59665f
C1434 dvdd.n51 dvss 1.29818f
C1435 dvdd.n52 dvss 1.40778f
C1436 dvdd.n53 dvss 0.046603f
C1437 dvdd.n54 dvss 0.046603f
C1438 dvdd.n55 dvss 2.85795f
C1439 dvdd.n56 dvss 2.85795f
C1440 dvdd.n57 dvss 0.043496f
C1441 dvdd.n58 dvss 0.043496f
C1442 dvdd.n59 dvss 0.043496f
C1443 dvdd.n60 dvss 0.04971f
C1444 dvdd.n61 dvss 0.04971f
C1445 dvdd.n64 dvss 0.04971f
C1446 dvdd.n68 dvss 0.030994f
C1447 dvdd.n69 dvss 0.030994f
C1448 dvdd.n70 dvss 1.6282f
C1449 dvdd.n71 dvss 0.043496f
C1450 dvdd.n72 dvss 0.043496f
C1451 dvdd.n73 dvss 0.043496f
C1452 dvdd.n74 dvss 0.027887f
C1453 dvdd.n79 dvss 0.286123f
C1454 dvdd.n89 dvss 0.043496f
C1455 dvdd.n93 dvss 0.030994f
C1456 dvdd.n94 dvss 0.030994f
C1457 dvdd.n96 dvss 0.04971f
C1458 dvdd.n97 dvss 1.6282f
C1459 dvdd.n98 dvss 0.043496f
C1460 dvdd.n99 dvss 0.043496f
C1461 dvdd.n100 dvss 0.043496f
C1462 dvdd.n101 dvss 0.027887f
C1463 dvdd.n103 dvss 0.107873f
C1464 dvdd.n105 dvss 0.286123f
C1465 dvdd.n111 dvss 0.030994f
C1466 dvdd.n116 dvss 0.056513f
C1467 dvdd.n117 dvss 0.103756f
C1468 dvdd.t5 dvss 0.588209f
C1469 dvdd.n126 dvss 0.010144f
C1470 dvdd.n129 dvss 0.021012f
C1471 dvdd.n132 dvss 0.021012f
C1472 dvdd.n133 dvss 0.023532f
C1473 dvdd.n134 dvss 1.43542f
C1474 dvdd.n135 dvss 1.43542f
C1475 dvdd.n136 dvss 0.023532f
C1476 dvdd.n137 dvss 0.023532f
C1477 dvdd.n138 dvss 0.023532f
C1478 dvdd.n139 dvss 0.023532f
C1479 dvdd.n140 dvss 0.023532f
C1480 dvdd.n141 dvss 0.017905f
C1481 dvdd.n142 dvss 0.017905f
C1482 dvdd.n143 dvss 0.017905f
C1483 dvdd.n144 dvss 0.021012f
C1484 dvdd.n147 dvss 0.021012f
C1485 dvdd.n151 dvss 0.021012f
C1486 dvdd.n154 dvss 0.422397f
C1487 dvdd.n166 dvss 0.023532f
C1488 dvdd.n167 dvss 0.021012f
C1489 dvdd.n169 dvss 0.021012f
C1490 dvdd.n170 dvss 0.017905f
C1491 dvdd.n179 dvss 0.156383f
C1492 dvdd.n182 dvss 0.021012f
C1493 dvdd.n185 dvss 0.021012f
C1494 dvdd.n187 dvss 0.023532f
C1495 dvdd.n188 dvss 0.021012f
C1496 dvdd.n191 dvss 0.021012f
C1497 dvdd.n193 dvss 0.017905f
C1498 dvdd.n195 dvss 0.010144f
C1499 dvdd.n196 dvss 0.017905f
C1500 dvdd.n197 dvss 0.023532f
C1501 dvdd.n198 dvss 0.017905f
C1502 dvdd.n201 dvss 0.021012f
C1503 dvdd.n204 dvss 0.021012f
C1504 dvdd.n216 dvss 0.021012f
C1505 dvdd.n219 dvss 0.023532f
C1506 dvdd.n220 dvss 0.021012f
C1507 dvdd.t37 dvss 0.588209f
C1508 dvdd.n227 dvss 0.021012f
C1509 dvdd.n230 dvss 0.021012f
C1510 dvdd.n231 dvss 0.023532f
C1511 dvdd.n232 dvss 0.021012f
C1512 dvdd.n236 dvss 0.021012f
C1513 dvdd.n239 dvss 0.017905f
C1514 dvdd.n240 dvss 0.023532f
C1515 dvdd.n241 dvss 0.023532f
C1516 dvdd.t1 dvss 2.28264f
C1517 dvdd.n242 dvss 0.023532f
C1518 dvdd.n243 dvss 0.021012f
C1519 dvdd.n247 dvss 0.100936f
C1520 dvdd.n248 dvss 0.103756f
C1521 dvdd.n249 dvss 0.100936f
C1522 dvdd.n250 dvss 0.103756f
C1523 dvdd.n251 dvss 0.100936f
C1524 dvdd.n252 dvss 0.110606f
C1525 dvdd.n253 dvss 0.156383f
C1526 dvdd.n255 dvss 0.422397f
C1527 dvdd.n257 dvss 0.09771f
C1528 dvdd.n258 dvss 0.053786f
C1529 dvdd.n260 dvss 0.032678f
C1530 dvdd.n261 dvss 0.016786f
C1531 dvdd.n262 dvss 0.017819f
C1532 dvdd.n263 dvss 0.017819f
C1533 dvdd.n264 dvss 0.119483f
C1534 dvdd.n265 dvss 0.060247f
C1535 dvdd.n267 dvss 0.074464f
C1536 dvdd.t116 dvss 0.452132f
C1537 dvdd.n268 dvss 0.270747f
C1538 dvdd.n269 dvss 0.032678f
C1539 dvdd.n270 dvss 0.322893f
C1540 dvdd.n271 dvss 0.093187f
C1541 dvdd.n273 dvss 0.074464f
C1542 dvdd.t106 dvss 0.218923f
C1543 dvdd.n274 dvss 0.140612f
C1544 dvdd.n275 dvss 0.028056f
C1545 dvdd.n276 dvss 0.203261f
C1546 dvdd.n277 dvss 0.0328f
C1547 dvdd.n278 dvss 0.010645f
C1548 dvdd.n279 dvss 0.0328f
C1549 dvdd.n280 dvss 0.036043f
C1550 dvdd.n281 dvss 0.015273f
C1551 dvdd.n282 dvss 0.032851f
C1552 dvdd.n283 dvss 0.010645f
C1553 dvdd.n284 dvss 0.010645f
C1554 dvdd.n285 dvss 0.014705f
C1555 dvdd.n286 dvss 0.010645f
C1556 dvdd.n289 dvss 0.014317f
C1557 dvdd.n290 dvss 0.011074f
C1558 dvdd.n291 dvss 0.010645f
C1559 dvdd.n292 dvss 0.010645f
C1560 dvdd.n294 dvss 0.010645f
C1561 dvdd.n295 dvss 0.010645f
C1562 dvdd.n296 dvss 0.029238f
C1563 dvdd.n297 dvss 0.033729f
C1564 dvdd.n299 dvss 0.010645f
C1565 dvdd.n301 dvss 0.010645f
C1566 dvdd.n303 dvss 0.010645f
C1567 dvdd.n305 dvss 0.010645f
C1568 dvdd.n307 dvss 0.010645f
C1569 dvdd.n309 dvss 0.010645f
C1570 dvdd.n311 dvss 0.010645f
C1571 dvdd.n313 dvss 0.010645f
C1572 dvdd.n315 dvss 0.014317f
C1573 dvdd.n318 dvss 0.010645f
C1574 dvdd.n319 dvss 0.010645f
C1575 dvdd.n320 dvss 0.023922f
C1576 dvdd.n321 dvss 0.018042f
C1577 dvdd.n322 dvss 0.020224f
C1578 dvdd.n323 dvss 0.010645f
C1579 dvdd.n324 dvss 0.010645f
C1580 dvdd.n325 dvss 0.014705f
C1581 dvdd.n326 dvss 0.010645f
C1582 dvdd.t47 dvss 0.047118f
C1583 dvdd.n328 dvss 0.017491f
C1584 dvdd.n329 dvss 0.013193f
C1585 dvdd.n332 dvss 0.010645f
C1586 dvdd.n334 dvss 0.010645f
C1587 dvdd.n336 dvss 0.010645f
C1588 dvdd.n338 dvss 0.010645f
C1589 dvdd.n340 dvss 0.010645f
C1590 dvdd.n342 dvss 0.010645f
C1591 dvdd.n344 dvss 0.010645f
C1592 dvdd.n346 dvss 0.010645f
C1593 dvdd.n347 dvss 0.014705f
C1594 dvdd.n348 dvss 0.010645f
C1595 dvdd.n349 dvss 0.023862f
C1596 dvdd.n351 dvss 0.013193f
C1597 dvdd.t36 dvss 0.047118f
C1598 dvdd.n352 dvss 0.017491f
C1599 dvdd.n354 dvss 0.020224f
C1600 dvdd.n355 dvss 0.017921f
C1601 dvdd.n356 dvss 0.023862f
C1602 dvdd.n357 dvss 0.12185f
C1603 dvdd.t89 dvss 0.354048f
C1604 dvdd.n358 dvss 0.12185f
C1605 dvdd.n359 dvss 0.020224f
C1606 dvdd.n360 dvss 0.011074f
C1607 dvdd.n362 dvss 0.014705f
C1608 dvdd.t62 dvss 0.047118f
C1609 dvdd.n363 dvss 0.014705f
C1610 dvdd.n366 dvss 0.014705f
C1611 dvdd.t68 dvss 0.047118f
C1612 dvdd.n367 dvss 0.014705f
C1613 dvdd.n370 dvss 0.014705f
C1614 dvdd.t86 dvss 0.047118f
C1615 dvdd.n371 dvss 0.014705f
C1616 dvdd.n374 dvss 0.014705f
C1617 dvdd.t40 dvss 0.047118f
C1618 dvdd.n375 dvss 0.014705f
C1619 dvdd.n377 dvss 0.011074f
C1620 dvdd.n378 dvss 0.020224f
C1621 dvdd.n379 dvss 0.121833f
C1622 dvdd.t0 dvss 0.354048f
C1623 dvdd.n380 dvss 0.121833f
C1624 dvdd.n381 dvss 0.023922f
C1625 dvdd.n383 dvss 0.010645f
C1626 dvdd.n385 dvss 0.010645f
C1627 dvdd.t100 dvss 0.02469f
C1628 dvdd.n386 dvss 0.111795f
C1629 dvdd.t33 dvss 0.047118f
C1630 dvdd.n388 dvss 0.014705f
C1631 dvdd.n389 dvss 0.017134f
C1632 dvdd.n390 dvss 0.017134f
C1633 dvdd.n391 dvss 0.014705f
C1634 dvdd.t83 dvss 0.047118f
C1635 dvdd.n392 dvss 0.014705f
C1636 dvdd.t80 dvss 0.047118f
C1637 dvdd.n395 dvss 0.014705f
C1638 dvdd.n397 dvss 0.010645f
C1639 dvdd.n398 dvss 0.010645f
C1640 dvdd.n399 dvss 0.075221f
C1641 dvdd.n400 dvss 0.075221f
C1642 dvdd.n402 dvss 0.014317f
C1643 dvdd.t11 dvss 0.047118f
C1644 dvdd.n403 dvss 0.014705f
C1645 dvdd.n406 dvss 0.014705f
C1646 dvdd.t8 dvss 0.047118f
C1647 dvdd.n407 dvss 0.014705f
C1648 dvdd.n410 dvss 0.014705f
C1649 dvdd.t4 dvss 0.047118f
C1650 dvdd.n411 dvss 0.014705f
C1651 dvdd.n414 dvss 0.014705f
C1652 dvdd.t77 dvss 0.047118f
C1653 dvdd.n415 dvss 0.014705f
C1654 dvdd.n417 dvss 0.065873f
C1655 dvdd.n418 dvss 0.037022f
C1656 dvdd.n419 dvss 0.071883f
C1657 dvdd.n420 dvss 0.375183f
C1658 dvdd.n421 dvss 1.52361f
C1659 dvdd.n422 dvss 0.081677f
C1660 dvdd.n423 dvss 0.308032f
C1661 dvdd.n424 dvss 12.7602f
C1662 dvdd.n425 dvss 1.35293f
C1663 dvdd.n427 dvss 0.013575f
C1664 dvdd.n428 dvss 0.010645f
C1665 dvdd.n429 dvss 0.036043f
C1666 dvdd.n430 dvss 0.041463f
C1667 dvdd.n431 dvss 0.014615f
C1668 dvdd.n432 dvss 0.042441f
C1669 dvdd.n433 dvss 0.010645f
C1670 dvdd.n435 dvss 0.010645f
C1671 dvdd.n436 dvss 0.015273f
C1672 dvdd.n437 dvss 0.010645f
C1673 dvdd.n438 dvss 0.0328f
C1674 dvdd.n439 dvss 0.036043f
C1675 dvdd.n440 dvss 0.244097f
C1676 dvdd.t65 dvss 0.705513f
C1677 dvdd.n441 dvss 0.2444f
C1678 dvdd.n442 dvss 0.036043f
C1679 dvdd.n443 dvss 0.010146f
C1680 dvdd.n444 dvss 0.010645f
C1681 dvdd.n446 dvss 0.010645f
C1682 dvdd.n448 dvss 0.010645f
C1683 dvdd.n450 dvss 0.010645f
C1684 dvdd.n452 dvss 0.013193f
C1685 dvdd.n453 dvss 0.010146f
C1686 dvdd.n454 dvss 0.010645f
C1687 dvdd.n455 dvss 0.015273f
C1688 dvdd.n456 dvss 0.036043f
C1689 dvdd.n457 dvss 0.2444f
C1690 dvdd.t43 dvss 0.705513f
C1691 dvdd.n458 dvss 0.2444f
C1692 dvdd.n459 dvss 0.036043f
C1693 dvdd.n461 dvss 0.017491f
C1694 dvdd.t22 dvss 0.047118f
C1695 dvdd.n462 dvss 0.014705f
C1696 dvdd.n465 dvss 0.014705f
C1697 dvdd.t18 dvss 0.047118f
C1698 dvdd.n466 dvss 0.014705f
C1699 dvdd.n469 dvss 0.014705f
C1700 dvdd.t71 dvss 0.047118f
C1701 dvdd.n470 dvss 0.014705f
C1702 dvdd.n473 dvss 0.014705f
C1703 dvdd.t53 dvss 0.047118f
C1704 dvdd.n474 dvss 0.014705f
C1705 dvdd.n476 dvss 0.223971f
C1706 dvdd.n477 dvss 0.081677f
C1707 dvdd.n478 dvss 1.49529f
C1708 dvdd.n479 dvss 1.27502f
C1709 dvdd.n480 dvss 0.045334f
C1710 dvdd.n481 dvss 0.244249f
C1711 dvdd.t56 dvss 0.705513f
C1712 dvdd.n482 dvss 0.2444f
C1713 dvdd.n483 dvss 0.035514f
C1714 dvdd.n484 dvss 0.035924f
C1715 dvdd.n485 dvss 0.248685f
C1716 dvdd.t50 dvss 0.705513f
C1717 dvdd.n486 dvss 0.2444f
C1718 dvdd.n487 dvss 0.033729f
C1719 dvdd.n489 dvss 0.014705f
C1720 dvdd.t59 dvss 0.047118f
C1721 dvdd.n490 dvss 0.014705f
C1722 dvdd.t74 dvss 0.047118f
C1723 dvdd.n493 dvss 0.014705f
C1724 dvdd.n495 dvss 0.010645f
C1725 dvdd.n498 dvss 0.014317f
C1726 dvdd.t29 dvss 0.047118f
C1727 dvdd.n499 dvss 0.014705f
C1728 dvdd.n501 dvss 0.011074f
C1729 dvdd.n502 dvss 0.033729f
C1730 dvdd.n503 dvss 0.2444f
C1731 dvdd.t14 dvss 0.705513f
C1732 dvdd.n504 dvss 0.225848f
C1733 dvdd.n505 dvss 0.090993f
C1734 dvdd.n506 dvss 0.024986f
C1735 dvdd.n507 dvss 0.065326f
C1736 dvdd.n508 dvss 0.091048f
C1737 dvdd.n509 dvss 0.022671f
C1738 dvdd.n510 dvss 0.010645f
C1739 dvdd.n511 dvss 0.0328f
C1740 dvdd.t25 dvss 0.705513f
C1741 dvdd.n512 dvss 0.2444f
C1742 dvdd.n513 dvss 0.036043f
C1743 dvdd.n514 dvss 0.015273f
C1744 dvdd.n515 dvss 0.027822f
C1745 dvdd.n516 dvss 0.049973f
C1746 dvdd.n517 dvss 0.064787f
C1747 dvdd.n518 dvss 0.143915f
C1748 dvdd.n519 dvss 0.140612f
C1749 dvdd.n520 dvss 0.014162f
C1750 dvdd.n521 dvss 0.207443f
C1751 dvdd.n522 dvss 0.014162f
C1752 dvdd.n523 dvss 0.168738f
C1753 dvdd.n527 dvss 0.04971f
C1754 dvdd.n528 dvss 0.046603f
C1755 dvdd.n533 dvss 0.030994f
C1756 dvdd.n534 dvss 0.027887f
C1757 dvdd.n537 dvss 0.030994f
C1758 dvdd.n538 dvss 0.043496f
C1759 dvdd.n539 dvss 0.04971f
C1760 dvdd.n540 dvss 0.043496f
C1761 dvdd.n541 dvss 0.04971f
C1762 dvdd.n543 dvss 0.04971f
C1763 dvdd.n545 dvss 0.04971f
C1764 dvdd.n546 dvss 0.046603f
C1765 dvdd.n550 dvss 0.027887f
C1766 dvdd.n551 dvss 0.043496f
C1767 dvdd.n552 dvss 0.039337f
C1768 dvdd.n553 dvss 0.107355f
C1769 dvdd.n554 dvss 0.140612f
C1770 dvdd.n555 dvss 0.113454f
C1771 dvdd.n556 dvss 0.036594f
C1772 dvdd.n557 dvss 0.06246f
C1773 dvdd.t108 dvss 0.900486f
C1774 dvdd.n559 dvss 0.61011f
C1775 dvdd.n560 dvss 0.06246f
C1776 dvdd.n562 dvss 0.61011f
C1777 dvdd.n563 dvss 0.028056f
C1778 dvdd.n564 dvss 0.037624f
C1779 dvdd.n565 dvss 0.19485f
C1780 dvdd.n566 dvss 0.127092f
C1781 dvdd.n567 dvss 0.014314f
C1782 dvdd.t94 dvss 0.213183f
C1783 dvdd.n569 dvss 0.014314f
C1784 dvdd.n570 dvss 0.07779f
C1785 dvdd.n571 dvss 0.064054f
C1786 dvdd.n572 dvss 0.122394f
C1787 dvdd.n573 dvss 0.154134f
C1788 dvdd.n574 dvss 0.014314f
C1789 dvdd.t119 dvss 0.213183f
C1790 dvdd.n576 dvss 0.014314f
C1791 dvdd.n577 dvss 0.142335f
C1792 dvdd.n578 dvss 0.080996f
C1793 dvdd.n579 dvss 0.050207f
C1794 dvdd.n580 dvss 0.010631f
C1795 dvdd.n581 dvss 0.017574f
C1796 dvdd.n583 dvss 0.140612f
C1797 dvdd.n584 dvss 0.017574f
C1798 dvdd.n585 dvss 0.137506f
C1799 dvdd.n586 dvss 0.240599f
C1800 dvdd.n587 dvss 0.162376f
C1801 dvdd.n588 dvss 0.181751f
C1802 dvdd.n589 dvss 0.029923f
C1803 dvdd.n591 dvss 0.270747f
C1804 dvdd.n592 dvss 0.029923f
C1805 dvdd.n593 dvss 0.023108f
C1806 dvdd.n594 dvss 0.037797f
C1807 dvdd.n595 dvss 0.049199f
C1808 dvdd.n596 dvss 0.141164f
C1809 dvdd.t99 dvss 0.203824f
C1810 dvdd.n599 dvss 0.141164f
C1811 dvdd.n600 dvss 0.016845f
C1812 dvdd.n601 dvss 0.046178f
C1813 dvdd.n613 dvss 0.043496f
C1814 dvdd.n614 dvss 0.030994f
C1815 dvdd.t30 dvss 0.398441f
C1816 dvdd.n618 dvss 0.195832f
C1817 dvdd.n619 dvss 0.803358f
C1818 dvdd.n620 dvss 1.40467f
C1819 dvdd.n621 dvss 0.043496f
C1820 dvdd.t15 dvss 2.85795f
C1821 dvdd.n622 dvss 0.043496f
C1822 dvdd.n623 dvss 0.043496f
C1823 dvdd.n624 dvss 0.04971f
C1824 dvdd.n625 dvss 0.043496f
C1825 dvdd.n626 dvss 0.04971f
C1826 dvdd.n627 dvss 0.043496f
C1827 dvdd.n629 dvss 0.030994f
C1828 dvdd.n632 dvss 0.030994f
C1829 dvdd.n633 dvss 0.027887f
C1830 dvdd.n635 dvss 0.030994f
C1831 dvdd.n638 dvss 0.030994f
C1832 dvdd.t19 dvss 0.398441f
C1833 dvdd.n650 dvss 0.30719f
C1834 dvdd.n651 dvss 0.803358f
C1835 dvdd.n652 dvss 1.40467f
C1836 dvdd.n653 dvss 0.043496f
C1837 dvdd.t44 dvss 2.85795f
C1838 dvdd.n654 dvss 0.043496f
C1839 dvdd.n655 dvss 0.043496f
C1840 dvdd.n656 dvss 0.04971f
C1841 dvdd.n657 dvss 0.043496f
C1842 dvdd.n658 dvss 0.043496f
C1843 dvdd.t26 dvss 2.85795f
C1844 dvdd.n659 dvss 0.043496f
C1845 dvdd.n660 dvss 0.811936f
C1846 dvdd.n661 dvss 0.702335f
C1847 dvdd.n662 dvss 3.31573f
C1848 dvdd.n663 dvss 14.948f
C1849 dvdd.n664 dvss 5.33263f
C1850 dvdd.n665 dvss 2.76314f
C1851 dvdd.n666 dvss 0.967096f
C1852 dvdd.n667 dvss 1.10126f
C1853 multiplexer_0.vtrip_1_b.n0 dvss 1.52802f
C1854 multiplexer_0.vtrip_1_b.t0 dvss 0.083414f
C1855 multiplexer_0.vtrip_1_b.t1 dvss 0.043789f
C1856 multiplexer_0.vtrip_1_b.t4 dvss 0.05762f
C1857 multiplexer_0.vtrip_1_b.t10 dvss 0.727869f
C1858 multiplexer_0.vtrip_1_b.t9 dvss 0.756194f
C1859 multiplexer_0.vtrip_1_b.t2 dvss 0.056412f
C1860 multiplexer_0.vtrip_1_b.t11 dvss 0.727869f
C1861 multiplexer_0.vtrip_1_b.t8 dvss 0.756194f
C1862 multiplexer_0.vtrip_1_b.t7 dvss 0.727869f
C1863 multiplexer_0.vtrip_1_b.t5 dvss 0.756194f
C1864 multiplexer_0.vtrip_1_b.t3 dvss 0.727869f
C1865 multiplexer_0.vtrip_1_b.t12 dvss 0.756194f
C1866 multiplexer_0.vtrip_1_b.t6 dvss 0.758654f
C1867 avss.t75 dvss 0.107061f
C1868 avss.n0 dvss 1.30263f
C1869 avss.t122 dvss 0.107275f
C1870 avss.t48 dvss 0.107061f
C1871 avss.t28 dvss 0.107061f
C1872 avss.t253 dvss 0.107061f
C1873 avss.t38 dvss 0.107061f
C1874 avss.t11 dvss 0.107061f
C1875 avss.t210 dvss 0.107061f
C1876 avss.t137 dvss 0.107061f
C1877 avss.t204 dvss 0.107061f
C1878 avss.t60 dvss 0.107061f
C1879 avss.t248 dvss 0.107061f
C1880 avss.t70 dvss 0.107061f
C1881 avss.t230 dvss 0.107061f
C1882 avss.t124 dvss 0.107061f
C1883 avss.t63 dvss 0.107061f
C1884 avss.t212 dvss 0.107061f
C1885 avss.t228 dvss 0.107061f
C1886 avss.t101 dvss 0.107061f
C1887 avss.t115 dvss 0.107061f
C1888 avss.t236 dvss 0.107061f
C1889 avss.t126 dvss 0.107061f
C1890 avss.t200 dvss 0.107061f
C1891 avss.t135 dvss 0.107061f
C1892 avss.t157 dvss 0.107061f
C1893 avss.t170 dvss 0.107061f
C1894 avss.t143 dvss 0.107061f
C1895 avss.t208 dvss 0.107061f
C1896 avss.t177 dvss 0.107061f
C1897 avss.t79 dvss 0.107061f
C1898 avss.t93 dvss 0.107061f
C1899 avss.t111 dvss 0.107061f
C1900 avss.t119 dvss 0.107061f
C1901 avss.t206 dvss 0.107061f
C1902 avss.t4 dvss 0.107061f
C1903 avss.t105 dvss 0.107061f
C1904 avss.t145 dvss 0.107061f
C1905 avss.t73 dvss 0.107061f
C1906 avss.t181 dvss 0.107061f
C1907 avss.t139 dvss 0.107061f
C1908 avss.t36 dvss 0.107061f
C1909 avss.t14 dvss 0.107061f
C1910 avss.t40 dvss 0.107061f
C1911 avss.t255 dvss 0.107061f
C1912 avss.t183 dvss 0.107061f
C1913 avss.t165 dvss 0.107061f
C1914 avss.t215 dvss 0.107061f
C1915 avss.t91 dvss 0.107061f
C1916 avss.t196 dvss 0.118399f
C1917 avss.t88 dvss 0.107275f
C1918 avss.n1 dvss 1.88827f
C1919 avss.t87 dvss 0.107061f
C1920 avss.n2 dvss 1.88849f
C1921 avss.t197 dvss 0.107275f
C1922 avss.n3 dvss 0.841011f
C1923 avss.n4 dvss 1.38053f
C1924 avss.t92 dvss 0.107275f
C1925 avss.n5 dvss 1.9273f
C1926 avss.t216 dvss 0.107275f
C1927 avss.n6 dvss 2.12999f
C1928 avss.t166 dvss 0.107275f
C1929 avss.n7 dvss 2.12999f
C1930 avss.t184 dvss 0.107275f
C1931 avss.n8 dvss 2.12999f
C1932 avss.t256 dvss 0.107275f
C1933 avss.n9 dvss 2.12999f
C1934 avss.t41 dvss 0.107275f
C1935 avss.n10 dvss 2.12999f
C1936 avss.t15 dvss 0.107275f
C1937 avss.n11 dvss 2.12999f
C1938 avss.t37 dvss 0.107275f
C1939 avss.n12 dvss 2.12999f
C1940 avss.t140 dvss 0.107275f
C1941 avss.n13 dvss 2.12999f
C1942 avss.t182 dvss 0.107275f
C1943 avss.n14 dvss 2.12999f
C1944 avss.t74 dvss 0.107275f
C1945 avss.n15 dvss 2.12999f
C1946 avss.t146 dvss 0.107275f
C1947 avss.n16 dvss 2.12999f
C1948 avss.t106 dvss 0.107275f
C1949 avss.n17 dvss 2.12999f
C1950 avss.t5 dvss 0.107275f
C1951 avss.n18 dvss 2.12999f
C1952 avss.t207 dvss 0.107275f
C1953 avss.n19 dvss 2.12999f
C1954 avss.t120 dvss 0.107275f
C1955 avss.n20 dvss 2.12999f
C1956 avss.t112 dvss 0.107275f
C1957 avss.n21 dvss 2.12999f
C1958 avss.t94 dvss 0.107275f
C1959 avss.n22 dvss 2.12999f
C1960 avss.t80 dvss 0.107275f
C1961 avss.n23 dvss 2.12999f
C1962 avss.t178 dvss 0.107275f
C1963 avss.n24 dvss 2.12999f
C1964 avss.t209 dvss 0.107275f
C1965 avss.n25 dvss 2.12999f
C1966 avss.t144 dvss 0.107275f
C1967 avss.n26 dvss 2.12999f
C1968 avss.t171 dvss 0.107275f
C1969 avss.n27 dvss 2.12999f
C1970 avss.t158 dvss 0.107275f
C1971 avss.n28 dvss 2.12999f
C1972 avss.t136 dvss 0.107275f
C1973 avss.n29 dvss 2.12999f
C1974 avss.t201 dvss 0.107275f
C1975 avss.n30 dvss 2.12999f
C1976 avss.t127 dvss 0.107275f
C1977 avss.n31 dvss 2.12999f
C1978 avss.t237 dvss 0.107275f
C1979 avss.n32 dvss 2.12999f
C1980 avss.t116 dvss 0.107275f
C1981 avss.n33 dvss 2.12999f
C1982 avss.t102 dvss 0.107275f
C1983 avss.n34 dvss 2.12999f
C1984 avss.t229 dvss 0.107275f
C1985 avss.n35 dvss 2.12999f
C1986 avss.t213 dvss 0.107275f
C1987 avss.n36 dvss 2.12999f
C1988 avss.t64 dvss 0.107275f
C1989 avss.n37 dvss 2.12999f
C1990 avss.t125 dvss 0.107275f
C1991 avss.n38 dvss 2.12999f
C1992 avss.t231 dvss 0.107275f
C1993 avss.n39 dvss 2.12999f
C1994 avss.t71 dvss 0.107275f
C1995 avss.n40 dvss 2.12999f
C1996 avss.t249 dvss 0.107275f
C1997 avss.n41 dvss 2.12999f
C1998 avss.t61 dvss 0.107275f
C1999 avss.n42 dvss 2.12999f
C2000 avss.t205 dvss 0.107275f
C2001 avss.n43 dvss 2.12999f
C2002 avss.t138 dvss 0.107275f
C2003 avss.n44 dvss 2.12999f
C2004 avss.t211 dvss 0.107275f
C2005 avss.n45 dvss 2.12999f
C2006 avss.t12 dvss 0.107275f
C2007 avss.n46 dvss 2.12999f
C2008 avss.t39 dvss 0.107275f
C2009 avss.n47 dvss 2.12999f
C2010 avss.t254 dvss 0.107275f
C2011 avss.n48 dvss 2.12999f
C2012 avss.t29 dvss 0.107275f
C2013 avss.n49 dvss 2.12999f
C2014 avss.t49 dvss 0.107275f
C2015 avss.n50 dvss 2.12999f
C2016 avss.t121 dvss 0.107061f
C2017 avss.n51 dvss 2.10879f
C2018 avss.t133 dvss 0.107061f
C2019 avss.n52 dvss 1.80989f
C2020 avss.t134 dvss 0.107275f
C2021 avss.n53 dvss 1.88827f
C2022 avss.t65 dvss 0.107061f
C2023 avss.n54 dvss 1.88849f
C2024 avss.t66 dvss 0.107275f
C2025 avss.n55 dvss 1.88827f
C2026 avss.t217 dvss 0.107061f
C2027 avss.n56 dvss 1.88849f
C2028 avss.t218 dvss 0.107275f
C2029 avss.n57 dvss 1.80931f
C2030 avss.t198 dvss 0.107061f
C2031 avss.t199 dvss 0.107275f
C2032 avss.n58 dvss 2.10843f
C2033 avss.t44 dvss 0.107061f
C2034 avss.t45 dvss 0.107275f
C2035 avss.n59 dvss 2.12999f
C2036 avss.t241 dvss 0.107061f
C2037 avss.t242 dvss 0.107275f
C2038 avss.n60 dvss 2.12999f
C2039 avss.t52 dvss 0.107061f
C2040 avss.t53 dvss 0.107275f
C2041 avss.n61 dvss 2.12999f
C2042 avss.t251 dvss 0.107061f
C2043 avss.t252 dvss 0.107275f
C2044 avss.n62 dvss 2.12999f
C2045 avss.t30 dvss 0.107061f
C2046 avss.t31 dvss 0.107275f
C2047 avss.n63 dvss 2.12999f
C2048 avss.t50 dvss 0.107061f
C2049 avss.t51 dvss 0.107275f
C2050 avss.n64 dvss 2.12999f
C2051 avss.t172 dvss 0.107061f
C2052 avss.t173 dvss 0.107275f
C2053 avss.n65 dvss 2.12999f
C2054 avss.t151 dvss 0.107061f
C2055 avss.t152 dvss 0.107275f
C2056 avss.n66 dvss 2.12999f
C2057 avss.t9 dvss 0.107061f
C2058 avss.t10 dvss 0.107275f
C2059 avss.n67 dvss 2.12999f
C2060 avss.t77 dvss 0.107061f
C2061 avss.t78 dvss 0.107275f
C2062 avss.n68 dvss 2.12999f
C2063 avss.t57 dvss 0.107061f
C2064 avss.t58 dvss 0.107275f
C2065 avss.n69 dvss 2.12999f
C2066 avss.t220 dvss 0.107061f
C2067 avss.t221 dvss 0.107275f
C2068 avss.n70 dvss 2.12999f
C2069 avss.t34 dvss 0.107061f
C2070 avss.t35 dvss 0.107275f
C2071 avss.n71 dvss 2.12999f
C2072 avss.t148 dvss 0.107061f
C2073 avss.t149 dvss 0.107275f
C2074 avss.n72 dvss 2.12999f
C2075 avss.t85 dvss 0.107061f
C2076 avss.t86 dvss 0.107275f
C2077 avss.n73 dvss 2.12999f
C2078 avss.t159 dvss 0.107061f
C2079 avss.t160 dvss 0.107275f
C2080 avss.n74 dvss 2.12999f
C2081 avss.t67 dvss 0.107061f
C2082 avss.t68 dvss 0.107275f
C2083 avss.n75 dvss 2.12999f
C2084 avss.t81 dvss 0.107061f
C2085 avss.t82 dvss 0.107275f
C2086 avss.n76 dvss 2.12999f
C2087 avss.t225 dvss 0.107061f
C2088 avss.t226 dvss 0.107275f
C2089 avss.n77 dvss 2.12999f
C2090 avss.t113 dvss 0.107061f
C2091 avss.t114 dvss 0.107275f
C2092 avss.n78 dvss 2.12999f
C2093 avss.t117 dvss 0.107061f
C2094 avss.t118 dvss 0.107275f
C2095 avss.n79 dvss 2.12999f
C2096 avss.t245 dvss 0.107061f
C2097 avss.t246 dvss 0.107275f
C2098 avss.n80 dvss 2.12999f
C2099 avss.t192 dvss 0.107061f
C2100 avss.t193 dvss 0.107275f
C2101 avss.n81 dvss 2.12999f
C2102 avss.t154 dvss 0.107061f
C2103 avss.t155 dvss 0.107275f
C2104 avss.n82 dvss 2.12999f
C2105 avss.t46 dvss 0.107061f
C2106 avss.t47 dvss 0.107275f
C2107 avss.n83 dvss 2.12999f
C2108 avss.t32 dvss 0.107061f
C2109 avss.t33 dvss 0.107275f
C2110 avss.n84 dvss 2.12999f
C2111 avss.t190 dvss 0.107061f
C2112 avss.t191 dvss 0.107275f
C2113 avss.n85 dvss 2.12999f
C2114 avss.t42 dvss 0.107061f
C2115 avss.t43 dvss 0.107275f
C2116 avss.n86 dvss 2.12999f
C2117 avss.t243 dvss 0.107061f
C2118 avss.t244 dvss 0.107275f
C2119 avss.n87 dvss 2.12999f
C2120 avss.t232 dvss 0.107061f
C2121 avss.t233 dvss 0.107275f
C2122 avss.n88 dvss 2.12999f
C2123 avss.t179 dvss 0.107061f
C2124 avss.t180 dvss 0.107275f
C2125 avss.n89 dvss 2.12999f
C2126 avss.t141 dvss 0.107061f
C2127 avss.t142 dvss 0.107275f
C2128 avss.n90 dvss 2.12999f
C2129 avss.t163 dvss 0.107061f
C2130 avss.t164 dvss 0.107275f
C2131 avss.n91 dvss 2.12999f
C2132 avss.t202 dvss 0.107061f
C2133 avss.t203 dvss 0.107275f
C2134 avss.n92 dvss 2.12999f
C2135 avss.t26 dvss 0.107061f
C2136 avss.t27 dvss 0.107275f
C2137 avss.n93 dvss 2.12999f
C2138 avss.t96 dvss 0.107061f
C2139 avss.t97 dvss 0.107275f
C2140 avss.n94 dvss 2.12999f
C2141 avss.t21 dvss 0.107061f
C2142 avss.t22 dvss 0.107275f
C2143 avss.n95 dvss 2.12999f
C2144 avss.t54 dvss 0.107061f
C2145 avss.t55 dvss 0.107275f
C2146 avss.n96 dvss 2.12999f
C2147 avss.t194 dvss 0.107061f
C2148 avss.t195 dvss 0.107275f
C2149 avss.n97 dvss 2.12999f
C2150 avss.t234 dvss 0.107061f
C2151 avss.t235 dvss 0.107275f
C2152 avss.n98 dvss 2.12999f
C2153 avss.t103 dvss 0.107061f
C2154 avss.t104 dvss 0.107275f
C2155 avss.n99 dvss 2.12999f
C2156 avss.t89 dvss 0.107061f
C2157 avss.t90 dvss 0.107275f
C2158 avss.n100 dvss 2.12999f
C2159 avss.t257 dvss 0.107061f
C2160 avss.t258 dvss 0.107275f
C2161 avss.n101 dvss 2.12999f
C2162 avss.t83 dvss 0.107061f
C2163 avss.t84 dvss 0.107275f
C2164 avss.n102 dvss 2.12999f
C2165 avss.t174 dvss 0.107061f
C2166 avss.t175 dvss 0.107275f
C2167 avss.n103 dvss 2.12999f
C2168 avss.t17 dvss 0.107061f
C2169 avss.t18 dvss 0.107275f
C2170 avss.n104 dvss 1.9273f
C2171 avss.t110 dvss 0.118589f
C2172 avss.n105 dvss 1.37998f
C2173 avss.t109 dvss 0.107061f
C2174 avss.n106 dvss 0.840861f
C2175 avss.t239 dvss 0.107275f
C2176 avss.n107 dvss 1.88827f
C2177 avss.t238 dvss 0.107061f
C2178 avss.n108 dvss 1.88849f
C2179 avss.t76 dvss 0.107275f
C2180 avss.n109 dvss 1.30278f
C2181 avss.n110 dvss 37.6986f
C2182 avss.n111 dvss 9.978429f
C2183 avss.n112 dvss 6.26811f
C2184 avss.n113 dvss 2.40542f
C2185 avss.n114 dvss 58.557697f
C2186 avss.t8 dvss 37.5956f
C2187 avss.t0 dvss 86.8916f
C2188 avss.n115 dvss 0.246751f
C2189 avss.n116 dvss 0.270556f
C2190 avss.n117 dvss 0.143093f
C2191 avss.n118 dvss 0.143093f
C2192 avss.n119 dvss 15.6291f
C2193 avss.t1 dvss 86.8916f
C2194 avss.t3 dvss 47.4543f
C2195 avss.n120 dvss 21.4327f
C2196 avss.n121 dvss 15.521199f
C2197 avss.n122 dvss 0.166279f
C2198 avss.n123 dvss 0.113061f
C2199 avss.t224 dvss 0.085003f
C2200 avss.n124 dvss 0.579451f
C2201 avss.n125 dvss 0.620407f
C2202 avss.n126 dvss 0.672677f
C2203 avss.n127 dvss 0.913668f
C2204 avss.n128 dvss 1.12574f
C2205 avss.t72 dvss 0.05686f
C2206 avss.t240 dvss 0.052438f
C2207 avss.n129 dvss 0.584392f
C2208 avss.n130 dvss 0.280151f
C2209 avss.n131 dvss 0.054797f
C2210 avss.n132 dvss 0.093477f
C2211 avss.n133 dvss 0.127609f
C2212 avss.t6 dvss 5.01586f
C2213 avss.n134 dvss 0.091567f
C2214 avss.n135 dvss 0.091567f
C2215 avss.n136 dvss 0.091567f
C2216 avss.n137 dvss 6.15944f
C2217 avss.n138 dvss 0.091567f
C2218 avss.n139 dvss 0.091567f
C2219 avss.n140 dvss 0.091567f
C2220 avss.n141 dvss 0.127609f
C2221 avss.n142 dvss 0.093477f
C2222 avss.n143 dvss 0.485764f
C2223 avss.n144 dvss 0.040626f
C2224 avss.n145 dvss 0.280151f
C2225 avss.t25 dvss 0.05686f
C2226 avss.t222 dvss 0.052438f
C2227 avss.n146 dvss 0.584392f
C2228 avss.t169 dvss 0.05686f
C2229 avss.t69 dvss 0.052438f
C2230 avss.n147 dvss 0.584392f
C2231 avss.n148 dvss 0.280151f
C2232 avss.n149 dvss 0.058072f
C2233 avss.n150 dvss 0.054797f
C2234 avss.n151 dvss 0.127609f
C2235 avss.n152 dvss 0.058265f
C2236 avss.n153 dvss 0.091567f
C2237 avss.n154 dvss 0.127609f
C2238 avss.n155 dvss 0.485764f
C2239 avss.n156 dvss 0.058072f
C2240 avss.n157 dvss 0.127609f
C2241 avss.n158 dvss 0.091567f
C2242 avss.n159 dvss 0.091567f
C2243 avss.n160 dvss 0.091567f
C2244 avss.n161 dvss 18.7238f
C2245 avss.n162 dvss 9.93295f
C2246 avss.t227 dvss 3.84753f
C2247 avss.n163 dvss 0.111972f
C2248 avss.n164 dvss 0.111972f
C2249 avss.n165 dvss 0.061622f
C2250 avss.n166 dvss 0.333049f
C2251 avss.n167 dvss 2.75401f
C2252 avss.t250 dvss 0.264743f
C2253 avss.n168 dvss 3.27009f
C2254 avss.n169 dvss 0.395908f
C2255 avss.n170 dvss 0.384325f
C2256 avss.n171 dvss 0.011407f
C2257 avss.n172 dvss 0.019304f
C2258 avss.n173 dvss 0.018536f
C2259 avss.n174 dvss 0.018536f
C2260 avss.n175 dvss 0.018536f
C2261 avss.n176 dvss 0.010661f
C2262 avss.n177 dvss 0.019304f
C2263 avss.n178 dvss 0.018536f
C2264 avss.n179 dvss 0.025823f
C2265 avss.n180 dvss 0.019304f
C2266 avss.n181 dvss 0.025052f
C2267 avss.n183 dvss 0.3173f
C2268 avss.n184 dvss 0.042212f
C2269 avss.n185 dvss 0.25032f
C2270 avss.n186 dvss 0.061622f
C2271 avss.n187 dvss 0.110471f
C2272 avss.n188 dvss 0.111972f
C2273 avss.n189 dvss 0.067664f
C2274 avss.n190 dvss 0.114349f
C2275 avss.n191 dvss 0.325415f
C2276 avss.t13 dvss 0.152677f
C2277 avss.t214 dvss 0.975027f
C2278 avss.n192 dvss 0.111972f
C2279 avss.n193 dvss 0.111972f
C2280 avss.n194 dvss 0.061622f
C2281 avss.n195 dvss 0.734956f
C2282 avss.n196 dvss 0.114349f
C2283 avss.n197 dvss 0.28176f
C2284 avss.n198 dvss 0.110471f
C2285 avss.n199 dvss 0.067664f
C2286 avss.n200 dvss 0.114349f
C2287 avss.n201 dvss 0.757068f
C2288 avss.n202 dvss 0.390643f
C2289 avss.t24 dvss 2.89879f
C2290 avss.n203 dvss 0.111972f
C2291 avss.n204 dvss 0.111972f
C2292 avss.n205 dvss 0.061622f
C2293 avss.n206 dvss 2.62332f
C2294 avss.n207 dvss 0.114349f
C2295 avss.n208 dvss 0.481981f
C2296 avss.n209 dvss 0.28176f
C2297 avss.n210 dvss 0.110471f
C2298 avss.n211 dvss 0.067664f
C2299 avss.n212 dvss 0.114349f
C2300 avss.n213 dvss 2.61079f
C2301 avss.n214 dvss 3.15651f
C2302 avss.t19 dvss 0.26454f
C2303 avss.n215 dvss 1.06406f
C2304 avss.t153 dvss 7.624569f
C2305 avss.n216 dvss 0.111972f
C2306 avss.n217 dvss 0.111972f
C2307 avss.n218 dvss 0.061622f
C2308 avss.n219 dvss 0.114349f
C2309 avss.n220 dvss 0.28176f
C2310 avss.n221 dvss 0.110471f
C2311 avss.n222 dvss 0.067664f
C2312 avss.n223 dvss 0.114349f
C2313 avss.n224 dvss 6.86705f
C2314 avss.n225 dvss 3.43526f
C2315 avss.t108 dvss 0.975027f
C2316 avss.n226 dvss 0.111972f
C2317 avss.n227 dvss 0.111972f
C2318 avss.n228 dvss 0.061622f
C2319 avss.n229 dvss 0.110471f
C2320 avss.n230 dvss 0.061622f
C2321 avss.n231 dvss 0.114349f
C2322 avss.n232 dvss 0.067664f
C2323 avss.n233 dvss 0.114349f
C2324 avss.n234 dvss 0.587544f
C2325 avss.n235 dvss 1.94342f
C2326 avss.n236 dvss 0.067664f
C2327 avss.n237 dvss 0.114349f
C2328 avss.n238 dvss 0.883421f
C2329 avss.n239 dvss 1.94342f
C2330 avss.t167 dvss 0.975027f
C2331 avss.n240 dvss 0.111972f
C2332 avss.n241 dvss 0.111972f
C2333 avss.n242 dvss 0.061622f
C2334 avss.n243 dvss 0.110471f
C2335 avss.n244 dvss 0.061622f
C2336 avss.n245 dvss 0.114349f
C2337 avss.n246 dvss 0.067664f
C2338 avss.n247 dvss 0.114349f
C2339 avss.n248 dvss 0.883421f
C2340 avss.n249 dvss 1.33105f
C2341 avss.n250 dvss 0.067664f
C2342 avss.n251 dvss 0.114349f
C2343 avss.n252 dvss 0.860256f
C2344 avss.n253 dvss 1.80693f
C2345 avss.t128 dvss 0.975027f
C2346 avss.n254 dvss 0.111972f
C2347 avss.n255 dvss 0.111972f
C2348 avss.n256 dvss 0.061622f
C2349 avss.n257 dvss 0.110471f
C2350 avss.n258 dvss 0.078068f
C2351 avss.n259 dvss 0.114349f
C2352 avss.n260 dvss 0.010661f
C2353 avss.n261 dvss 0.098021f
C2354 avss.n262 dvss 0.019304f
C2355 avss.n263 dvss 0.025052f
C2356 avss.t95 dvss 0.923456f
C2357 avss.n264 dvss 4.1063f
C2358 avss.n265 dvss 0.018536f
C2359 avss.n266 dvss 0.01795f
C2360 avss.n267 dvss 0.011407f
C2361 avss.n268 dvss 0.019304f
C2362 avss.t123 dvss 5.7008f
C2363 avss.n269 dvss 0.111972f
C2364 avss.n270 dvss 0.111972f
C2365 avss.n271 dvss 0.061622f
C2366 avss.n272 dvss 1.37613f
C2367 avss.n273 dvss 0.018536f
C2368 avss.n274 dvss 0.025052f
C2369 avss.n275 dvss 0.019304f
C2370 avss.n276 dvss 0.025856f
C2371 avss.n277 dvss 0.010661f
C2372 avss.n278 dvss 0.018536f
C2373 avss.n279 dvss 0.018536f
C2374 avss.t187 dvss 5.7008f
C2375 avss.n280 dvss 0.111972f
C2376 avss.n281 dvss 0.111972f
C2377 avss.n282 dvss 0.061622f
C2378 avss.n283 dvss 0.114349f
C2379 avss.n284 dvss 0.28176f
C2380 avss.n285 dvss 0.110471f
C2381 avss.n286 dvss 0.067664f
C2382 avss.n287 dvss 0.114349f
C2383 avss.n288 dvss 4.35256f
C2384 avss.n289 dvss 2.30248f
C2385 avss.n290 dvss 0.019304f
C2386 avss.n291 dvss 0.018536f
C2387 avss.n292 dvss 0.018536f
C2388 avss.n293 dvss 0.019304f
C2389 avss.n294 dvss 0.011407f
C2390 avss.t98 dvss 0.812642f
C2391 avss.n295 dvss 0.025052f
C2392 avss.n296 dvss 0.025856f
C2393 avss.n297 dvss 0.044004f
C2394 avss.n298 dvss 0.035359f
C2395 avss.n299 dvss 0.044004f
C2396 avss.n300 dvss 0.018536f
C2397 avss.n301 dvss 2.3148f
C2398 avss.n302 dvss 4.37718f
C2399 avss.n303 dvss 0.114349f
C2400 avss.n304 dvss 0.280952f
C2401 avss.n305 dvss 0.28176f
C2402 avss.n306 dvss 0.110471f
C2403 avss.n307 dvss 0.067664f
C2404 avss.n308 dvss 0.114349f
C2405 avss.n309 dvss 4.35256f
C2406 avss.n310 dvss 2.17936f
C2407 avss.n311 dvss 0.018536f
C2408 avss.n312 dvss 0.018536f
C2409 avss.n313 dvss 0.019304f
C2410 avss.n314 dvss 0.018536f
C2411 avss.n315 dvss 0.067664f
C2412 avss.n316 dvss 0.114349f
C2413 avss.n317 dvss 17.3824f
C2414 avss.n318 dvss 0.587544f
C2415 avss.n319 dvss 0.587544f
C2416 avss.n320 dvss 0.587544f
C2417 avss.n321 dvss 0.067664f
C2418 avss.n322 dvss 0.114349f
C2419 avss.n323 dvss 0.587544f
C2420 avss.n324 dvss 0.587544f
C2421 avss.n325 dvss 0.587544f
C2422 avss.t130 dvss 0.975027f
C2423 avss.n326 dvss 0.111972f
C2424 avss.n327 dvss 0.111972f
C2425 avss.n328 dvss 0.061622f
C2426 avss.n329 dvss 0.860256f
C2427 avss.n330 dvss 0.114349f
C2428 avss.n331 dvss 0.044004f
C2429 avss.n332 dvss 0.044004f
C2430 avss.n333 dvss 0.019304f
C2431 avss.n334 dvss 0.019304f
C2432 avss.n335 dvss 0.019304f
C2433 avss.n336 dvss 0.356546f
C2434 avss.n337 dvss 0.018536f
C2435 avss.n338 dvss 0.025052f
C2436 avss.n339 dvss 0.025856f
C2437 avss.n340 dvss 0.018536f
C2438 avss.n341 dvss 0.018536f
C2439 avss.n342 dvss 0.418019f
C2440 avss.n343 dvss 0.018536f
C2441 avss.n344 dvss 0.018536f
C2442 avss.n345 dvss 0.018536f
C2443 avss.n346 dvss 0.025856f
C2444 avss.n347 dvss 0.025052f
C2445 avss.t131 dvss 0.153684f
C2446 avss.n348 dvss 0.011407f
C2447 avss.n349 dvss 0.010661f
C2448 avss.n350 dvss 0.035359f
C2449 avss.n351 dvss 0.272575f
C2450 avss.n352 dvss 0.061622f
C2451 avss.n353 dvss 0.114349f
C2452 avss.n354 dvss 0.067664f
C2453 avss.n355 dvss 0.114349f
C2454 avss.n356 dvss 1.80693f
C2455 avss.t161 dvss 0.975027f
C2456 avss.n357 dvss 0.111972f
C2457 avss.n358 dvss 0.111972f
C2458 avss.n359 dvss 0.061622f
C2459 avss.n360 dvss 0.114349f
C2460 avss.n361 dvss 0.061622f
C2461 avss.n362 dvss 0.114349f
C2462 avss.n363 dvss 0.067664f
C2463 avss.n364 dvss 0.114349f
C2464 avss.t162 dvss 0.975027f
C2465 avss.n365 dvss 0.111972f
C2466 avss.n366 dvss 0.111972f
C2467 avss.n367 dvss 0.061622f
C2468 avss.n368 dvss 0.110471f
C2469 avss.n369 dvss 0.061622f
C2470 avss.n370 dvss 0.114349f
C2471 avss.n371 dvss 0.067664f
C2472 avss.n372 dvss 0.114349f
C2473 avss.n373 dvss 0.883421f
C2474 avss.n374 dvss 0.067664f
C2475 avss.n375 dvss 0.114349f
C2476 avss.n376 dvss 0.860256f
C2477 avss.n377 dvss 1.80693f
C2478 avss.t20 dvss 0.975027f
C2479 avss.n378 dvss 0.111972f
C2480 avss.n379 dvss 0.111972f
C2481 avss.n380 dvss 0.061622f
C2482 avss.n381 dvss 0.114349f
C2483 avss.n382 dvss 0.067664f
C2484 avss.n383 dvss 0.110471f
C2485 avss.n384 dvss 0.061622f
C2486 avss.n385 dvss 0.114349f
C2487 avss.n386 dvss 0.067664f
C2488 avss.n387 dvss 0.114349f
C2489 avss.n388 dvss 0.860256f
C2490 avss.n389 dvss 0.111972f
C2491 avss.t147 dvss 0.975027f
C2492 avss.n390 dvss 0.111972f
C2493 avss.n391 dvss 0.110471f
C2494 avss.n392 dvss 0.28176f
C2495 avss.n393 dvss 0.24099f
C2496 avss.n394 dvss 0.061622f
C2497 avss.n395 dvss 0.114349f
C2498 avss.n396 dvss 0.067664f
C2499 avss.n397 dvss 0.114349f
C2500 avss.n398 dvss 0.860256f
C2501 avss.n399 dvss 0.111972f
C2502 avss.t62 dvss 0.975027f
C2503 avss.n400 dvss 0.111972f
C2504 avss.n401 dvss 0.110471f
C2505 avss.n402 dvss 0.28176f
C2506 avss.n403 dvss 0.24099f
C2507 avss.n404 dvss 0.061622f
C2508 avss.n405 dvss 0.114349f
C2509 avss.n406 dvss 0.067664f
C2510 avss.n407 dvss 0.114349f
C2511 avss.n408 dvss 0.860256f
C2512 avss.n409 dvss 0.111972f
C2513 avss.t247 dvss 0.975027f
C2514 avss.n410 dvss 0.111972f
C2515 avss.n411 dvss 0.110471f
C2516 avss.n412 dvss 0.28176f
C2517 avss.n413 dvss 0.24099f
C2518 avss.n414 dvss 0.24099f
C2519 avss.n415 dvss 0.28176f
C2520 avss.n416 dvss 0.114349f
C2521 avss.n417 dvss 0.860256f
C2522 avss.n418 dvss 1.80693f
C2523 avss.n419 dvss 0.860256f
C2524 avss.n420 dvss 0.111972f
C2525 avss.t219 dvss 0.975027f
C2526 avss.n421 dvss 0.111972f
C2527 avss.n422 dvss 0.110471f
C2528 avss.n423 dvss 0.28176f
C2529 avss.n424 dvss 0.24099f
C2530 avss.n425 dvss 0.24099f
C2531 avss.n426 dvss 0.28176f
C2532 avss.n427 dvss 0.114349f
C2533 avss.n428 dvss 0.883421f
C2534 avss.n429 dvss 1.94342f
C2535 avss.n430 dvss 0.883421f
C2536 avss.n431 dvss 1.94342f
C2537 avss.t99 dvss 0.975027f
C2538 avss.n432 dvss 0.111972f
C2539 avss.n433 dvss 0.111972f
C2540 avss.n434 dvss 0.061622f
C2541 avss.n435 dvss 0.114349f
C2542 avss.n436 dvss 0.061622f
C2543 avss.n437 dvss 0.114349f
C2544 avss.n438 dvss 0.067664f
C2545 avss.n439 dvss 0.114349f
C2546 avss.n440 dvss 0.988598f
C2547 avss.t185 dvss 0.135242f
C2548 avss.n441 dvss 0.883421f
C2549 avss.n442 dvss 0.018536f
C2550 avss.n443 dvss 0.025052f
C2551 avss.n444 dvss 0.019304f
C2552 avss.n445 dvss 0.025856f
C2553 avss.n446 dvss 0.061622f
C2554 avss.n447 dvss 0.114349f
C2555 avss.n448 dvss 0.067664f
C2556 avss.n449 dvss 0.114349f
C2557 avss.n450 dvss 0.860256f
C2558 avss.n451 dvss 0.111972f
C2559 avss.t56 dvss 0.975027f
C2560 avss.n452 dvss 0.111972f
C2561 avss.n453 dvss 0.110471f
C2562 avss.n454 dvss 0.28176f
C2563 avss.n455 dvss 0.184828f
C2564 avss.n456 dvss 0.330663f
C2565 avss.n457 dvss 0.044004f
C2566 avss.n458 dvss 0.019304f
C2567 avss.n459 dvss 0.025052f
C2568 avss.n460 dvss 0.025856f
C2569 avss.n461 dvss 0.018536f
C2570 avss.n462 dvss 0.018536f
C2571 avss.n463 dvss 0.018536f
C2572 avss.n464 dvss 0.43851f
C2573 avss.n465 dvss 0.018536f
C2574 avss.n466 dvss 0.019304f
C2575 avss.n467 dvss 0.011407f
C2576 avss.n468 dvss 0.010661f
C2577 avss.n469 dvss 0.035359f
C2578 avss.n470 dvss 0.044004f
C2579 avss.n471 dvss 0.018536f
C2580 avss.n472 dvss 0.444658f
C2581 avss.t176 dvss 0.975027f
C2582 avss.n473 dvss 0.111972f
C2583 avss.n474 dvss 0.111972f
C2584 avss.n475 dvss 0.061622f
C2585 avss.n476 dvss 0.757068f
C2586 avss.n477 dvss 0.114349f
C2587 avss.n478 dvss 0.067664f
C2588 avss.n479 dvss 0.110471f
C2589 avss.n480 dvss 0.24099f
C2590 avss.n481 dvss 0.28176f
C2591 avss.n482 dvss 0.114349f
C2592 avss.n483 dvss 0.587544f
C2593 avss.n484 dvss 5.94779f
C2594 avss.n485 dvss 6.68171f
C2595 avss.n486 dvss 9.88291f
C2596 avss.n487 dvss 4.16193f
C2597 avss.n488 dvss 40.396103f
C2598 avss.n489 dvss 26.021599f
C2599 avss.n490 dvss 0.883421f
C2600 avss.n491 dvss 0.111972f
C2601 avss.t107 dvss 0.975027f
C2602 avss.n492 dvss 0.111972f
C2603 avss.n493 dvss 0.110471f
C2604 avss.n494 dvss 0.28176f
C2605 avss.n495 dvss 0.24099f
C2606 avss.n496 dvss 0.061622f
C2607 avss.n497 dvss 0.114349f
C2608 avss.n498 dvss 0.067664f
C2609 avss.n499 dvss 0.114349f
C2610 avss.n500 dvss 0.587544f
C2611 avss.n501 dvss 1.06406f
C2612 avss.n502 dvss 0.587544f
C2613 avss.n503 dvss 0.883421f
C2614 avss.n504 dvss 0.111972f
C2615 avss.t189 dvss 0.975027f
C2616 avss.n505 dvss 0.111972f
C2617 avss.n506 dvss 0.110471f
C2618 avss.n507 dvss 0.28176f
C2619 avss.n508 dvss 0.24099f
C2620 avss.n509 dvss 0.061622f
C2621 avss.n510 dvss 0.114349f
C2622 avss.n511 dvss 0.067664f
C2623 avss.n512 dvss 0.114349f
C2624 avss.n513 dvss 0.587544f
C2625 avss.n514 dvss 0.883421f
C2626 avss.n515 dvss 0.111972f
C2627 avss.t156 dvss 0.975027f
C2628 avss.n516 dvss 0.111972f
C2629 avss.n517 dvss 0.110471f
C2630 avss.n518 dvss 0.28176f
C2631 avss.n519 dvss 0.230303f
C2632 avss.n520 dvss 0.137752f
C2633 avss.n521 dvss 0.061622f
C2634 avss.n522 dvss 0.114349f
C2635 avss.n523 dvss 0.067664f
C2636 avss.n524 dvss 0.114349f
C2637 avss.n525 dvss 0.025052f
C2638 avss.n526 dvss 0.019304f
C2639 avss.n527 dvss 0.025714f
C2640 avss.n528 dvss 0.010661f
C2641 avss.n529 dvss 0.011407f
C2642 avss.n530 dvss 0.019304f
C2643 avss.n531 dvss 0.018536f
C2644 avss.n532 dvss 0.018536f
C2645 avss.n533 dvss 0.019304f
C2646 avss.n534 dvss 0.018536f
C2647 avss.n535 dvss 0.025714f
C2648 avss.n536 dvss 0.025052f
C2649 avss.n538 dvss 0.304183f
C2650 avss.n539 dvss 0.036852f
C2651 avss.n540 dvss 0.030559f
C2652 avss.n541 dvss 0.036852f
C2653 avss.n542 dvss 0.018536f
C2654 avss.n543 dvss 0.374849f
C2655 avss.n544 dvss 0.725479f
C2656 avss.n545 dvss 0.883421f
C2657 avss.n546 dvss 0.111972f
C2658 avss.t188 dvss 0.975027f
C2659 avss.n547 dvss 0.111972f
C2660 avss.n548 dvss 0.110471f
C2661 avss.n549 dvss 0.28176f
C2662 avss.n550 dvss 0.25032f
C2663 avss.n551 dvss 0.24099f
C2664 avss.n552 dvss 0.28176f
C2665 avss.n553 dvss 0.110471f
C2666 avss.n554 dvss 0.067664f
C2667 avss.n555 dvss 0.114349f
C2668 avss.n556 dvss 0.883421f
C2669 avss.n557 dvss 1.94342f
C2670 avss.n558 dvss 0.883421f
C2671 avss.n559 dvss 0.860256f
C2672 avss.n560 dvss 0.111972f
C2673 avss.t59 dvss 0.975027f
C2674 avss.n561 dvss 0.111972f
C2675 avss.n562 dvss 0.110471f
C2676 avss.n563 dvss 0.28176f
C2677 avss.n564 dvss 0.24099f
C2678 avss.n565 dvss 0.24099f
C2679 avss.n566 dvss 0.28176f
C2680 avss.n567 dvss 0.110471f
C2681 avss.n568 dvss 0.067664f
C2682 avss.n569 dvss 0.114349f
C2683 avss.n570 dvss 0.860256f
C2684 avss.n571 dvss 1.80693f
C2685 avss.n572 dvss 0.860256f
C2686 avss.n573 dvss 0.111972f
C2687 avss.t168 dvss 0.975027f
C2688 avss.n574 dvss 0.111972f
C2689 avss.n575 dvss 0.110471f
C2690 avss.n576 dvss 0.28176f
C2691 avss.n577 dvss 0.24099f
C2692 avss.n578 dvss 0.186634f
C2693 avss.n579 dvss 0.28176f
C2694 avss.n580 dvss 0.110471f
C2695 avss.n581 dvss 0.067664f
C2696 avss.n582 dvss 0.114349f
C2697 avss.n583 dvss 0.587544f
C2698 avss.t100 dvss 7.01827f
C2699 avss.n584 dvss 0.025052f
C2700 avss.n585 dvss 6.64036f
C2701 avss.n586 dvss 0.024963f
C2702 avss.n587 dvss 0.025052f
C2703 avss.n588 dvss 0.296155f
C2704 avss.n589 dvss 0.064234f
C2705 avss.n590 dvss 0.024963f
C2706 avss.n591 dvss 4.83181f
C2707 avss.n592 dvss 9.85383f
C2708 avss.n593 dvss 3.43526f
C2709 avss.n594 dvss 0.090028f
C2710 avss.n595 dvss 0.111972f
C2711 avss.t150 dvss 5.7008f
C2712 avss.n596 dvss 0.111972f
C2713 avss.n597 dvss 0.054886f
C2714 avss.n598 dvss 0.070963f
C2715 avss.n599 dvss 0.019536f
C2716 avss.n600 dvss 0.025052f
C2717 avss.n601 dvss 0.018536f
C2718 avss.n602 dvss 2.05623f
C2719 avss.n603 dvss 0.018536f
C2720 avss.n604 dvss 0.090326f
C2721 avss.n605 dvss 0.059153f
C2722 avss.n606 dvss 0.050002f
C2723 avss.n607 dvss 0.243047f
C2724 avss.n608 dvss 0.24099f
C2725 avss.n609 dvss 0.28176f
C2726 avss.n610 dvss 0.114349f
C2727 avss.n611 dvss 0.860256f
C2728 avss.n612 dvss 1.80693f
C2729 avss.n613 dvss 0.860256f
C2730 avss.n614 dvss 0.111972f
C2731 avss.t16 dvss 0.975027f
C2732 avss.n615 dvss 0.111972f
C2733 avss.n616 dvss 0.110471f
C2734 avss.n617 dvss 0.28176f
C2735 avss.n618 dvss 0.24099f
C2736 avss.n619 dvss 0.24099f
C2737 avss.n620 dvss 0.28176f
C2738 avss.n621 dvss 0.114349f
C2739 avss.n622 dvss 0.883421f
C2740 avss.n623 dvss 1.94342f
C2741 avss.n624 dvss 0.883421f
C2742 avss.n625 dvss 0.111972f
C2743 avss.t186 dvss 0.975027f
C2744 avss.n626 dvss 0.111972f
C2745 avss.n627 dvss 0.110471f
C2746 avss.n628 dvss 0.28176f
C2747 avss.n629 dvss 0.24099f
C2748 avss.n630 dvss 0.24099f
C2749 avss.n631 dvss 0.28176f
C2750 avss.n632 dvss 0.114349f
C2751 avss.n633 dvss 0.587544f
C2752 avss.n634 dvss 2.95743f
C2753 avss.n635 dvss 5.89287f
C2754 avss.n636 dvss 3.56744f
C2755 avss.n637 dvss 2.61079f
C2756 avss.t23 dvss 2.89879f
C2757 avss.n638 dvss 0.111972f
C2758 avss.n639 dvss 0.114349f
C2759 avss.n640 dvss 0.28176f
C2760 avss.n641 dvss 0.471293f
C2761 avss.n642 dvss 0.137752f
C2762 avss.n643 dvss 0.034156f
C2763 avss.n644 dvss 0.042212f
C2764 avss.n645 dvss 0.025823f
C2765 avss.n646 dvss 0.025052f
C2766 avss.t129 dvss 0.147412f
C2767 avss.n647 dvss 4.16246f
C2768 avss.n648 dvss 3.48605f
C2769 avss.n649 dvss 0.114349f
C2770 avss.n650 dvss 0.067664f
C2771 avss.n651 dvss 0.110471f
C2772 avss.n652 dvss 0.41942f
C2773 avss.n653 dvss 0.114349f
C2774 avss.n654 dvss 2.48054f
C2775 avss.n655 dvss 38.3628f
C2776 avss.n656 dvss 33.1972f
C2777 avss.n657 dvss 6.21863f
C2778 avss.n658 dvss 6.23994f
C2779 avss.n659 dvss 0.127609f
C2780 avss.n660 dvss 0.093477f
C2781 avss.n661 dvss 0.058072f
C2782 avss.n662 dvss 0.485764f
C2783 avss.n663 dvss 0.058265f
C2784 avss.n664 dvss 0.069303f
C2785 avss.n665 dvss 0.040626f
C2786 avss.n666 dvss 0.054797f
C2787 avss.n667 dvss 0.058072f
C2788 avss.n668 dvss 0.091567f
C2789 avss.n669 dvss 0.127609f
C2790 avss.n670 dvss 0.093477f
C2791 avss.n671 dvss 0.485764f
C2792 avss.n672 dvss 0.058265f
C2793 avss.n673 dvss 0.058072f
C2794 avss.n674 dvss 0.127609f
C2795 avss.n675 dvss 0.280151f
C2796 avss.t132 dvss 0.05686f
C2797 avss.t7 dvss 0.052438f
C2798 avss.n676 dvss 0.584392f
C2799 avss.n677 dvss 0.23107f
C2800 avss.n678 dvss 0.22828f
C2801 avss.n679 dvss 0.279644f
C2802 avss.n680 dvss 0.058173f
C2803 avss.n681 dvss 0.054797f
C2804 avss.n682 dvss 0.093477f
C2805 avss.n683 dvss 0.069303f
C2806 avss.n684 dvss 0.040626f
C2807 avss.n685 dvss 0.054797f
C2808 avss.n686 dvss 0.058072f
C2809 avss.n687 dvss 0.091567f
C2810 avss.n688 dvss 0.069303f
C2811 avss.n689 dvss 0.093477f
C2812 avss.n690 dvss 0.058265f
C2813 avss.n691 dvss 0.054797f
C2814 avss.n692 dvss 0.058072f
C2815 avss.n693 dvss 0.091567f
C2816 avss.n694 dvss 8.86258f
C2817 avss.n695 dvss 0.091567f
C2818 avss.n696 dvss 0.093477f
C2819 avss.n697 dvss 0.093477f
C2820 avss.n698 dvss 0.069303f
C2821 avss.n699 dvss 0.040626f
C2822 avss.n700 dvss 0.054797f
C2823 avss.n701 dvss 0.058173f
C2824 avss.n702 dvss 0.279644f
C2825 avss.n703 dvss 0.22828f
C2826 avss.n704 dvss 0.23107f
C2827 avss.n705 dvss 1.18122f
C2828 avss.n706 dvss 0.789556f
C2829 avss.n707 dvss 0.22828f
C2830 avss.n708 dvss 0.279644f
C2831 avss.n709 dvss 0.058173f
C2832 avss.n710 dvss 0.054797f
C2833 avss.n711 dvss 0.058072f
C2834 avss.n712 dvss 0.091567f
C2835 avss.n713 dvss 6.30083f
C2836 avss.n714 dvss 0.091567f
C2837 avss.n715 dvss 0.058173f
C2838 avss.n716 dvss 0.279644f
C2839 avss.n717 dvss 0.22828f
C2840 avss.n718 dvss 0.23107f
C2841 avss.n719 dvss 3.95622f
C2842 avss.n720 dvss 21.1607f
C2843 avss.n721 dvss 6.11833f
C2844 avss.n722 dvss 6.03898f
C2845 avss.n723 dvss 5.55681f
C2846 avss.n724 dvss 5.75446f
C2847 avss.n725 dvss 1.45429f
C2848 avss.n726 dvss 1.4843f
C2849 avss.n727 dvss 1.79671f
C2850 avss.n728 dvss 0.143102f
C2851 avss.t223 dvss 24.9958f
C2852 avss.n729 dvss 0.143102f
C2853 avss.n730 dvss 0.109155f
C2854 avss.n731 dvss 1.84429f
C2855 avss.n732 dvss 4.9089f
C2856 avss.n733 dvss 6.53045f
C2857 avss.n734 dvss 2.40661f
C2858 avss.t2 dvss 86.8916f
C2859 avss.n735 dvss 2.40661f
C2860 avss.n736 dvss 24.0401f
C2861 avss.n737 dvss 10.747499f
C2862 avss.n738 dvss 13.144401f
C2863 avss.n739 dvss 16.679f
C2864 avss.n740 dvss 18.5431f
C2865 multiplexer_0.trans_gate_m_31.out.t0 dvss 2.86063f
C2866 multiplexer_0.trans_gate_m_31.out.t1 dvss 0.035046f
C2867 multiplexer_0.trans_gate_m_31.out.t4 dvss 0.035046f
C2868 multiplexer_0.trans_gate_m_31.out.t2 dvss 0.03423f
C2869 multiplexer_0.trans_gate_m_31.out.t3 dvss 0.035046f
C2870 multiplexer_0.trans_gate_m_29.in.t3 dvss 2.86081f
C2871 multiplexer_0.trans_gate_m_29.in.t2 dvss 0.035001f
C2872 multiplexer_0.trans_gate_m_29.in.t4 dvss 0.035001f
C2873 multiplexer_0.trans_gate_m_29.in.t1 dvss 0.034185f
C2874 multiplexer_0.trans_gate_m_29.in.t0 dvss 0.035001f
C2875 multiplexer_0.trans_gate_m_19.ena dvss 8.89849f
C2876 multiplexer_0.trans_gate_m_31.ena_b dvss 9.161139f
C2877 multiplexer_0.vtrip_1.n0 dvss 2.03852f
C2878 multiplexer_0.vtrip_1.t6 dvss 1.0902f
C2879 multiplexer_0.vtrip_1.t9 dvss 0.070793f
C2880 multiplexer_0.vtrip_1.t0 dvss 0.964007f
C2881 multiplexer_0.vtrip_1.t7 dvss 1.00152f
C2882 multiplexer_0.vtrip_1.t4 dvss 1.05073f
C2883 multiplexer_0.vtrip_1.t2 dvss 0.070793f
C2884 multiplexer_0.vtrip_1.t8 dvss 0.964007f
C2885 multiplexer_0.vtrip_1.t5 dvss 1.00152f
C2886 multiplexer_0.vtrip_1.t3 dvss 0.964007f
C2887 multiplexer_0.vtrip_1.t1 dvss 1.00152f
C2888 level_shifter_1.out dvss 8.02274f
.ends


magic
tech sky130A
magscale 1 2
timestamp 1713218293
<< metal1 >>
rect 339 2485 571 2543
rect 281 2427 397 2485
rect 513 2427 687 2485
rect 281 2369 339 2427
rect 629 2369 803 2427
rect 223 2079 339 2369
rect 745 2311 861 2369
rect 803 2253 919 2311
rect 861 2195 977 2253
rect 919 2138 1035 2195
rect 919 2137 1093 2138
rect 281 2021 339 2079
rect 977 2022 1093 2137
rect 1325 2080 1441 2138
rect 1267 2022 1441 2080
rect 281 1905 397 2021
rect 1035 1964 1151 2022
rect 1209 1964 1325 2022
rect 1093 1906 1267 1964
rect 223 1847 571 1905
rect 1035 1848 1151 1906
rect 165 1731 629 1847
rect 1035 1790 1093 1848
rect 977 1732 1093 1790
rect 165 1615 687 1731
rect 919 1674 1035 1732
rect 919 1616 977 1674
rect 165 1557 629 1615
rect 223 1499 629 1557
rect 861 1558 977 1616
rect 861 1500 919 1558
rect 281 1441 571 1499
rect 803 1442 919 1500
rect 1383 1499 1441 2022
rect 513 1383 571 1441
rect 745 1384 861 1442
rect 1383 1441 1499 1499
rect 745 1383 803 1384
rect 513 1325 629 1383
rect 687 1326 803 1383
rect 1325 1383 1499 1441
rect 687 1325 745 1326
rect 571 1209 745 1325
rect 1325 1325 1557 1383
rect 1325 1209 1383 1325
rect 1499 1267 1557 1325
rect 1499 1209 1615 1267
rect 629 1093 745 1209
rect 1267 1093 1383 1209
rect 1557 1151 1615 1209
rect 1557 1093 1673 1151
rect 571 1035 803 1093
rect 1267 1035 1325 1093
rect 571 919 629 1035
rect 745 977 803 1035
rect 1209 977 1325 1035
rect 1615 977 1673 1093
rect 745 919 861 977
rect 1209 919 1267 977
rect 1615 919 1731 977
rect 513 861 629 919
rect 803 861 919 919
rect 513 687 571 861
rect 861 803 919 861
rect 1151 861 1267 919
rect 1151 803 1209 861
rect 861 745 977 803
rect 1093 745 1209 803
rect 1673 803 1731 919
rect 1673 745 1789 803
rect 919 687 1035 745
rect 1093 687 1151 745
rect 455 629 571 687
rect 397 571 513 629
rect 339 513 513 571
rect 977 571 1151 687
rect 1731 571 1789 745
rect 977 513 1209 571
rect 281 455 397 513
rect 223 397 339 455
rect 165 339 281 397
rect 455 339 513 513
rect 919 397 1035 513
rect 1093 454 1209 513
rect 861 339 1035 397
rect 165 281 223 339
rect 107 223 223 281
rect 397 281 513 339
rect 803 281 919 339
rect 107 165 165 223
rect 49 107 165 165
rect 397 107 455 281
rect 803 224 861 281
rect 745 166 861 224
rect 687 108 803 166
rect 977 108 1035 339
rect 1151 396 1209 454
rect 1731 397 1847 571
rect 1151 338 1267 396
rect 1209 280 1325 338
rect 1789 281 1847 397
rect 1267 222 1383 280
rect 1673 223 1847 281
rect 1441 222 1499 223
rect 1325 165 1499 222
rect 1673 165 1789 223
rect 1325 164 1731 165
rect 49 49 107 107
rect 339 49 455 107
rect 629 50 745 108
rect 919 50 1035 108
rect 1441 107 1731 164
rect -9 -9 397 49
rect 571 -66 687 50
rect 629 -124 745 -66
rect 919 -124 977 50
rect 1499 49 1615 107
rect 687 -182 803 -124
rect 745 -240 803 -182
rect 861 -182 977 -124
rect 861 -240 919 -182
rect 745 -298 919 -240
rect 803 -356 861 -298
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713122376
<< nwell >>
rect -18218 17203 -2751 17489
rect -18218 -3716 -17932 17203
rect -3037 14033 -2751 17203
rect 7842 14053 24020 14339
rect -3037 13747 6011 14033
rect -3037 13726 -2751 13747
rect 5725 9115 6011 13747
rect 7842 10246 8128 14053
rect 7842 9960 11647 10246
rect 5725 8829 10262 9115
rect 9976 -3716 10262 8829
rect 11361 -130 11647 9960
rect 23734 -130 24020 14053
rect 11361 -416 24020 -130
rect -18218 -4000 10262 -3716
rect -18218 -4002 10239 -4000
use comp_hyst  comp_hyst_0
timestamp 1713115829
transform 1 0 6715 0 1 11235
box 1667 -5363 16947 2564
use level_shifter  level_shifter_0
timestamp 1713121837
transform 1 0 6519 0 1 8816
box 1105 -2314 6378 -340
use level_shifter  level_shifter_1
timestamp 1713121837
transform 1 0 6519 0 1 6624
box 1105 -2314 6378 -340
use level_shifter  level_shifter_2
timestamp 1713121837
transform 1 0 6519 0 1 4432
box 1105 -2314 6378 -340
use level_shifter  level_shifter_4
timestamp 1713121837
transform 1 0 6519 0 1 2240
box 1105 -2314 6378 -340
use multiplexer  multiplexer_0
timestamp 1713115829
transform 1 0 -1139 0 1 -203
box -199 -135 8108 13095
use voltage_divider  voltage_divider_0
timestamp 1713115829
transform 1 0 -16349 0 1 -2158
box -1259 -1438 14153 19128
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713017665
<< pwell >>
rect -183 -208 183 208
<< psubdiff >>
rect -147 138 -51 172
rect 51 138 147 172
rect -147 76 -113 138
rect 113 76 147 138
rect -147 -138 -113 -76
rect 113 -138 147 -76
rect -147 -172 -51 -138
rect 51 -172 147 -138
<< psubdiffcont >>
rect -51 138 51 172
rect -147 -76 -113 76
rect 113 -76 147 76
rect -51 -172 51 -138
<< ndiode >>
rect -45 58 45 70
rect -45 -58 -33 58
rect 33 -58 45 58
rect -45 -70 45 -58
<< ndiodec >>
rect -33 -58 33 58
<< locali >>
rect -147 138 -51 172
rect 51 138 147 172
rect -147 76 -113 138
rect 113 76 147 138
rect -33 58 33 74
rect -33 -74 33 -58
rect -147 -138 -113 -76
rect 113 -138 147 -76
rect -147 -172 -51 -138
rect 51 -172 147 -138
<< viali >>
rect -33 -58 33 58
<< metal1 >>
rect -39 58 39 70
rect -39 -58 -33 58
rect 33 -58 39 58
rect -39 -70 39 -58
<< properties >>
string FIXED_BBOX -130 -155 130 155
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 0.45 l 0.7 area 315.0m peri 2.3 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713121837
<< locali >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 2319 -509 3279 -340
rect 5235 -369 6338 -340
rect 5235 -492 5456 -369
rect 6301 -492 6338 -369
rect 5235 -538 6338 -492
rect 5235 -1104 5418 -538
rect 5234 -1740 5418 -1226
rect 1183 -2314 2143 -1781
rect 5551 -2034 6338 -1774
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 5234 -2121 6338 -2034
rect 5234 -2244 5276 -2121
rect 6276 -2244 6338 -2121
rect 5234 -2314 6338 -2244
<< viali >>
rect 1223 -493 2106 -370
rect 5456 -492 6301 -369
rect 2357 -2286 3240 -2163
rect 5276 -2244 6276 -2121
<< metal1 >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 5418 -369 6338 -340
rect 5418 -492 5456 -369
rect 6301 -492 6338 -369
rect 5418 -538 6338 -492
rect 1183 -758 1325 -539
rect 1353 -710 1363 -658
rect 1963 -710 1973 -658
rect 2489 -670 2499 -618
rect 3099 -670 3109 -618
rect 1183 -959 1357 -758
rect 1969 -830 2494 -746
rect 1969 -887 2205 -830
rect 2345 -887 2494 -830
rect 1969 -958 2494 -887
rect 1183 -1362 1325 -959
rect 1353 -1058 1363 -1006
rect 1963 -1058 1973 -1006
rect 2489 -1167 2505 -1151
rect 3095 -1167 3105 -1151
rect 2489 -1219 2499 -1167
rect 3099 -1219 3105 -1167
rect 1353 -1314 1363 -1262
rect 1963 -1314 1973 -1262
rect 1183 -1562 1357 -1362
rect 1969 -1427 2461 -1362
rect 1969 -1484 1985 -1427
rect 2125 -1484 2461 -1427
rect 2489 -1457 2499 -1405
rect 3099 -1457 3105 -1405
rect 2489 -1473 2504 -1457
rect 3095 -1473 3105 -1457
rect 1969 -1562 2461 -1484
rect 2462 -1562 2493 -1505
rect 1353 -1662 1363 -1610
rect 1963 -1662 1973 -1610
rect 2271 -1905 2493 -1562
rect 2489 -1953 3109 -1937
rect 2489 -2005 2499 -1953
rect 3099 -2005 3109 -1953
rect 3137 -2115 3279 -718
rect 5418 -721 5540 -538
rect 5568 -673 5578 -621
rect 6178 -673 6188 -621
rect 5418 -921 5572 -721
rect 6184 -921 6338 -721
rect 5568 -1021 5578 -969
rect 6178 -1021 6185 -969
rect 6213 -1104 6338 -921
rect 5452 -1225 6338 -1104
rect 5452 -1226 6304 -1225
rect 5452 -1400 5543 -1226
rect 5571 -1352 5577 -1300
rect 6178 -1352 6188 -1300
rect 5571 -1368 6188 -1352
rect 5452 -1599 5520 -1400
rect 5572 -1599 5582 -1400
rect 5452 -1600 5571 -1599
rect 6184 -1600 6338 -1400
rect 5568 -1700 5578 -1648
rect 6179 -1700 6189 -1648
rect 5326 -1926 5336 -1848
rect 5476 -1926 5486 -1848
rect 6217 -2034 6338 -1600
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 5234 -2121 6338 -2034
rect 5234 -2244 5276 -2121
rect 6276 -2244 6338 -2121
rect 5234 -2313 6338 -2244
rect 5234 -2314 5551 -2313
<< via1 >>
rect 1363 -710 1963 -658
rect 2499 -670 3099 -618
rect 2205 -887 2345 -830
rect 1363 -1058 1963 -1006
rect 2499 -1219 3099 -1167
rect 1363 -1314 1963 -1262
rect 1985 -1484 2125 -1427
rect 2499 -1457 3099 -1405
rect 1363 -1662 1963 -1610
rect 2499 -2005 3099 -1953
rect 5578 -673 6178 -621
rect 5578 -1021 6178 -969
rect 5577 -1352 6178 -1300
rect 5520 -1599 5572 -1400
rect 5578 -1700 6179 -1648
rect 5336 -1926 5476 -1848
<< metal2 >>
rect 2499 -616 6178 -606
rect 2499 -618 5339 -616
rect 1363 -657 2135 -643
rect 1363 -658 1985 -657
rect 1963 -710 1985 -658
rect 1363 -714 1985 -710
rect 2125 -714 2135 -657
rect 3099 -670 5339 -618
rect 2499 -673 5339 -670
rect 5479 -621 6178 -616
rect 5479 -673 5578 -621
rect 2499 -683 6178 -673
rect 1363 -720 2135 -714
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -897 2355 -887
rect 5327 -969 6178 -959
rect 1363 -1006 2135 -996
rect 1963 -1058 1985 -1006
rect 1363 -1063 1985 -1058
rect 2125 -1063 2135 -1006
rect 5327 -1026 5337 -969
rect 5477 -1021 5578 -969
rect 5477 -1026 6178 -1021
rect 5327 -1036 6178 -1026
rect 1363 -1068 2135 -1063
rect 1363 -1073 2125 -1068
rect 2499 -1164 5487 -1157
rect 2499 -1167 5337 -1164
rect 3099 -1219 5337 -1167
rect 2499 -1221 5337 -1219
rect 5477 -1221 5487 -1164
rect 2499 -1229 5487 -1221
rect 1363 -1257 2355 -1247
rect 1363 -1262 2205 -1257
rect 1963 -1314 2205 -1262
rect 2345 -1314 2355 -1257
rect 1363 -1324 2355 -1314
rect 5327 -1294 6178 -1285
rect 5327 -1351 5337 -1294
rect 5477 -1300 6178 -1294
rect 5477 -1351 5577 -1300
rect 5327 -1352 5577 -1351
rect 5327 -1362 6178 -1352
rect 2499 -1400 5572 -1390
rect 2499 -1405 3177 -1400
rect 1975 -1427 2135 -1417
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 3099 -1457 3177 -1405
rect 3317 -1457 5520 -1400
rect 2499 -1467 5520 -1457
rect 1975 -1494 2135 -1484
rect 1363 -1610 2355 -1600
rect 5520 -1609 5572 -1599
rect 1963 -1662 2205 -1610
rect 1363 -1667 2205 -1662
rect 2345 -1667 2355 -1610
rect 1363 -1672 2355 -1667
rect 5327 -1648 6179 -1638
rect 5327 -1705 5337 -1648
rect 5477 -1700 5578 -1648
rect 5477 -1705 6179 -1700
rect 5327 -1715 6179 -1705
rect 5336 -1848 5476 -1838
rect 5336 -1936 5476 -1926
rect 2499 -1952 3327 -1943
rect 2499 -1953 3177 -1952
rect 3099 -2005 3177 -1953
rect 2499 -2009 3177 -2005
rect 3317 -2009 3327 -1952
rect 2499 -2015 3327 -2009
<< via2 >>
rect 1985 -714 2125 -657
rect 5339 -673 5479 -616
rect 2205 -887 2345 -830
rect 1985 -1063 2125 -1006
rect 5337 -1026 5477 -969
rect 5337 -1221 5477 -1164
rect 2205 -1314 2345 -1257
rect 5337 -1351 5477 -1294
rect 1985 -1484 2125 -1427
rect 3177 -1457 3317 -1400
rect 2205 -1667 2345 -1610
rect 5337 -1705 5477 -1648
rect 5336 -1926 5476 -1848
rect 3177 -2009 3317 -1952
<< metal3 >>
rect 5327 -616 5488 -606
rect 1975 -657 2135 -648
rect 1975 -714 1985 -657
rect 2125 -714 2135 -657
rect 1975 -1006 2135 -714
rect 5327 -673 5339 -616
rect 5479 -673 5488 -616
rect 1975 -1063 1985 -1006
rect 2125 -1063 2135 -1006
rect 1975 -1427 2135 -1063
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 1975 -1494 2135 -1484
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -1257 2355 -887
rect 2195 -1314 2205 -1257
rect 2345 -1314 2355 -1257
rect 2195 -1610 2355 -1314
rect 5327 -969 5488 -673
rect 5327 -1026 5337 -969
rect 5477 -1026 5488 -969
rect 5327 -1164 5488 -1026
rect 5327 -1221 5337 -1164
rect 5477 -1221 5488 -1164
rect 5327 -1294 5488 -1221
rect 5327 -1351 5337 -1294
rect 5477 -1351 5488 -1294
rect 2195 -1667 2205 -1610
rect 2345 -1667 2355 -1610
rect 2195 -1672 2355 -1667
rect 3167 -1400 3327 -1390
rect 3167 -1457 3177 -1400
rect 3317 -1457 3327 -1400
rect 3167 -1952 3327 -1457
rect 5327 -1648 5488 -1351
rect 5327 -1705 5337 -1648
rect 5477 -1705 5488 -1648
rect 5327 -1843 5488 -1705
rect 5326 -1848 5488 -1843
rect 5326 -1926 5336 -1848
rect 5476 -1926 5488 -1848
rect 5326 -1931 5488 -1926
rect 3167 -2009 3177 -1952
rect 3317 -2009 3327 -1952
rect 3167 -2014 3327 -2009
rect 5327 -2015 5488 -1931
use sky130_fd_pr__diode_pw2nd_05v5_37RBXE  sky130_fd_pr__diode_pw2nd_05v5_37RBXE_0
timestamp 1713020003
transform 0 1 5406 -1 0 -1887
box -183 -208 183 208
use sky130_fd_pr__nfet_01v8_MG6U6H  sky130_fd_pr__nfet_01v8_MG6U6H_0
timestamp 1713020003
transform 1 0 5878 0 1 -1500
box -496 -310 496 310
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0
timestamp 1713020003
transform -1 0 2799 0 1 -1705
box -528 -458 528 458
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1
timestamp 1713020003
transform -1 0 2799 0 1 -919
box -528 -458 528 458
use sky130_fd_pr__pfet_01v8_J2L9Q3  sky130_fd_pr__pfet_01v8_J2L9Q3_0
timestamp 1713020003
transform 1 0 5878 0 1 -821
box -496 -319 496 319
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0
timestamp 1713020003
transform 1 0 1663 0 -1 -1462
box -558 -397 558 397
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1
timestamp 1713020003
transform 1 0 1663 0 -1 -858
box -558 -397 558 397
<< labels >>
flabel space 1105 -1255 2221 -461 0 FreeSans 1600 0 0 0 M3
flabel space 2271 -1377 3327 -461 0 FreeSans 1600 0 0 0 M5
flabel space 2271 -2163 3327 -1247 0 FreeSans 1600 0 0 0 M6
flabel metal1 1183 -539 2143 -340 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 1363 -1662 1963 -1610 0 FreeSans 800 0 0 0 out_b
port 2 nsew
flabel metal2 1363 -710 1963 -658 0 FreeSans 800 0 0 0 out
port 3 nsew
flabel space 1105 -1859 2221 -1065 0 FreeSans 1600 0 0 0 M4
flabel metal2 3317 -1467 3773 -1390 0 FreeSans 800 0 0 0 in_b
flabel metal1 2319 -2314 3279 -2115 0 FreeSans 1600 0 0 0 avss
port 4 nsew
flabel space 5418 -538 6378 -340 0 FreeSans 1600 0 0 0 dvdd
port 5 nsew
flabel metal3 5327 -2015 5488 -1926 0 FreeSans 1600 0 0 0 in
port 6 nsew
flabel space 5382 -1810 6374 -1190 0 FreeSans 1600 0 0 0 M1
flabel space 5382 -1140 6374 -502 0 FreeSans 1600 0 0 0 M2
flabel metal1 5234 -2313 6338 -2244 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
<< end >>

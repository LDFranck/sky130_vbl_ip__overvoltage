magic
tech sky130A
magscale 1 2
timestamp 1713147273
<< nwell >>
rect -18218 17203 -2751 17489
rect -18218 -3716 -17932 17203
rect -3037 14033 -2751 17203
rect 7842 14053 24078 14339
rect -3037 13747 6011 14033
rect 5725 9115 6011 13747
rect 7842 10246 8128 14053
rect 7842 9960 11647 10246
rect 5725 8829 10262 9115
rect 9976 -3716 10262 8829
rect 11361 -130 11647 9960
rect 23792 -130 24078 14053
rect 11361 -416 24078 -130
rect -18218 -4002 10262 -3716
<< nsubdiff >>
rect -18182 17433 -2831 17453
rect -18182 17399 -18100 17433
rect -2910 17399 -2831 17433
rect -18182 17379 -2831 17399
rect -18182 17373 -18108 17379
rect -18182 -3883 -18162 17373
rect -18128 -3883 -18108 17373
rect -2905 17358 -2831 17379
rect -2905 14008 -2885 17358
rect -2851 14008 -2831 17358
rect -2905 13997 -2831 14008
rect 7927 14283 24011 14303
rect 7927 14249 8003 14283
rect 23934 14249 24011 14283
rect 7927 14229 24011 14249
rect 7927 14223 8001 14229
rect -2905 13977 5975 13997
rect -2905 13943 -2831 13977
rect 5895 13943 5975 13977
rect -2905 13923 5975 13943
rect 5901 13919 5975 13923
rect 5901 9087 5921 13919
rect 5955 9087 5975 13919
rect 7927 10076 7947 14223
rect 7981 10076 8001 14223
rect 7927 10070 8001 10076
rect 23937 14223 24011 14229
rect 7927 10050 11472 10070
rect 7927 10016 8004 10050
rect 11396 10016 11472 10050
rect 7927 9996 11472 10016
rect 5901 9079 5975 9087
rect 11398 9990 11472 9996
rect 5901 9059 10225 9079
rect 5901 9025 5976 9059
rect 10148 9025 10225 9059
rect 5901 9005 10225 9025
rect -18182 -3891 -18108 -3883
rect 10151 8999 10225 9005
rect 10151 -3885 10171 8999
rect 10205 -3885 10225 8999
rect 11398 -299 11418 9990
rect 11452 -299 11472 9990
rect 11398 -305 11472 -299
rect 23937 -297 23957 14223
rect 23991 -297 24011 14223
rect 23937 -305 24011 -297
rect 11398 -325 24011 -305
rect 11398 -359 11478 -325
rect 23937 -359 24011 -325
rect 11398 -379 24011 -359
rect 10151 -3891 10225 -3885
rect -18182 -3912 10225 -3891
rect -18182 -3946 -18108 -3912
rect 10145 -3946 10225 -3912
rect -18182 -3965 10225 -3946
rect -18182 -3966 10217 -3965
<< nsubdiffcont >>
rect -18100 17399 -2910 17433
rect -18162 -3883 -18128 17373
rect -2885 14008 -2851 17358
rect 8003 14249 23934 14283
rect -2831 13943 5895 13977
rect 5921 9087 5955 13919
rect 7947 10076 7981 14223
rect 8004 10016 11396 10050
rect 5976 9025 10148 9059
rect 10171 -3885 10205 8999
rect 11418 -299 11452 9990
rect 23957 -297 23991 14223
rect 11478 -359 23937 -325
rect -18108 -3946 10145 -3912
<< locali >>
rect -18162 17399 -18100 17433
rect -2910 17399 -2851 17433
rect -18162 17373 -18128 17399
rect -2885 17358 -2851 17399
rect -2885 13977 -2851 14008
rect 7947 14249 8003 14283
rect 23934 14249 23991 14283
rect 7947 14223 7981 14249
rect -2885 13943 -2831 13977
rect 5895 13943 5955 13977
rect 5921 13919 5955 13943
rect 7947 10050 7981 10076
rect 23957 14223 23991 14249
rect 7947 10016 8004 10050
rect 11396 10016 11452 10050
rect 5921 9059 5955 9087
rect 11418 9990 11452 10016
rect 5921 9025 5976 9059
rect 10148 9025 10205 9059
rect -18162 -3912 -18128 -3883
rect 10171 8999 10205 9025
rect 11418 -325 11452 -299
rect 23957 -325 23991 -297
rect 11418 -359 11478 -325
rect 23937 -359 23991 -325
rect 10171 -3912 10205 -3885
rect -18162 -3946 -18108 -3912
rect 10145 -3945 10205 -3912
rect 10145 -3946 10204 -3945
<< metal2 >>
rect 2247 9698 7379 9775
rect 2215 9231 6918 9308
rect 7362 8170 7882 8173
rect 7362 8163 7892 8170
rect 7502 8106 7892 8163
rect 7362 8099 7892 8106
rect 7362 8096 7882 8099
<< via2 >>
rect 7362 8106 7502 8163
<< metal3 >>
rect 7352 8163 7512 8168
rect 7352 8106 7362 8163
rect 7502 8106 7512 8163
rect 7352 8101 7512 8106
use comp_hyst  comp_hyst_0
timestamp 1713115829
transform 1 0 6716 0 1 11234
box 1667 -5363 16947 2564
use level_shifter  level_shifter_0
timestamp 1713121837
transform 1 0 6519 0 1 8816
box 1105 -2314 6378 -340
use level_shifter  level_shifter_1
timestamp 1713121837
transform 1 0 6519 0 1 6624
box 1105 -2314 6378 -340
use level_shifter  level_shifter_2
timestamp 1713121837
transform 1 0 6519 0 1 4432
box 1105 -2314 6378 -340
use level_shifter  level_shifter_4
timestamp 1713121837
transform 1 0 6519 0 1 2240
box 1105 -2314 6378 -340
use multiplexer  multiplexer_0
timestamp 1713137003
transform 1 0 -1955 0 1 209
box -199 -135 8108 13095
use vd2mux_conn  vd2mux_conn_1
timestamp 1713130350
transform 1 0 478 0 1 1
box -3578 973 -2488 12383
use voltage_divider  voltage_divider_0
timestamp 1713115829
transform 1 0 -16053 0 1 -2158
box -1259 -1438 14153 19128
<< end >>

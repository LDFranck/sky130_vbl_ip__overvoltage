magic
tech sky130A
magscale 1 2
timestamp 1713017665
<< nwell >>
rect -1796 -319 1796 319
<< pmos >>
rect -1600 -100 1600 100
<< pdiff >>
rect -1658 88 -1600 100
rect -1658 -88 -1646 88
rect -1612 -88 -1600 88
rect -1658 -100 -1600 -88
rect 1600 88 1658 100
rect 1600 -88 1612 88
rect 1646 -88 1658 88
rect 1600 -100 1658 -88
<< pdiffc >>
rect -1646 -88 -1612 88
rect 1612 -88 1646 88
<< nsubdiff >>
rect -1760 249 -1664 283
rect 1664 249 1760 283
rect -1760 187 -1726 249
rect 1726 187 1760 249
rect -1760 -249 -1726 -187
rect 1726 -249 1760 -187
rect -1760 -283 -1664 -249
rect 1664 -283 1760 -249
<< nsubdiffcont >>
rect -1664 249 1664 283
rect -1760 -187 -1726 187
rect 1726 -187 1760 187
rect -1664 -283 1664 -249
<< poly >>
rect -1600 181 1600 197
rect -1600 147 -1584 181
rect 1584 147 1600 181
rect -1600 100 1600 147
rect -1600 -147 1600 -100
rect -1600 -181 -1584 -147
rect 1584 -181 1600 -147
rect -1600 -197 1600 -181
<< polycont >>
rect -1584 147 1584 181
rect -1584 -181 1584 -147
<< locali >>
rect -1760 249 -1664 283
rect 1664 249 1760 283
rect -1760 187 -1726 249
rect 1726 187 1760 249
rect -1600 147 -1584 181
rect 1584 147 1600 181
rect -1646 88 -1612 104
rect -1646 -104 -1612 -88
rect 1612 88 1646 104
rect 1612 -104 1646 -88
rect -1600 -181 -1584 -147
rect 1584 -181 1600 -147
rect -1760 -249 -1726 -187
rect 1726 -249 1760 -187
rect -1760 -283 -1664 -249
rect 1664 -283 1760 -249
<< viali >>
rect -1584 147 1584 181
rect -1646 -88 -1612 88
rect 1612 -88 1646 88
rect -1584 -181 1584 -147
<< metal1 >>
rect -1596 181 1596 187
rect -1596 147 -1584 181
rect 1584 147 1596 181
rect -1596 141 1596 147
rect -1652 88 -1606 100
rect -1652 -88 -1646 88
rect -1612 -88 -1606 88
rect -1652 -100 -1606 -88
rect 1606 88 1652 100
rect 1606 -88 1612 88
rect 1646 -88 1652 88
rect 1606 -100 1652 -88
rect -1596 -147 1596 -141
rect -1596 -181 -1584 -147
rect 1584 -181 1596 -147
rect -1596 -187 1596 -181
<< properties >>
string FIXED_BBOX -1743 -266 1743 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 16 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

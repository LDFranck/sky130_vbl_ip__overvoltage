magic
tech sky130A
magscale 1 2
timestamp 1713022109
<< locali >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 2319 -509 3279 -340
rect 3488 -369 4591 -340
rect 3488 -492 3709 -369
rect 4554 -492 4591 -369
rect 3488 -538 4591 -492
rect 3488 -1104 3671 -538
rect 3487 -1740 3671 -1226
rect 1183 -2314 2143 -1781
rect 3804 -2034 4591 -1774
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 3487 -2121 4591 -2034
rect 3487 -2244 3529 -2121
rect 4529 -2244 4591 -2121
rect 3487 -2314 4591 -2244
<< viali >>
rect 1223 -493 2106 -370
rect 3709 -492 4554 -369
rect 2357 -2286 3240 -2163
rect 3529 -2244 4529 -2121
<< metal1 >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 3671 -369 4591 -340
rect 3671 -492 3709 -369
rect 4554 -492 4591 -369
rect 3671 -538 4591 -492
rect 1183 -758 1325 -539
rect 1353 -710 1363 -658
rect 1963 -710 1973 -658
rect 2489 -670 2499 -618
rect 3099 -670 3109 -618
rect 1183 -959 1357 -758
rect 1969 -830 2494 -746
rect 1969 -887 2205 -830
rect 2345 -887 2494 -830
rect 1969 -958 2494 -887
rect 1183 -1362 1325 -959
rect 1353 -1058 1363 -1006
rect 1963 -1058 1973 -1006
rect 2489 -1167 2505 -1151
rect 3095 -1167 3105 -1151
rect 2489 -1219 2499 -1167
rect 3099 -1219 3105 -1167
rect 1353 -1314 1363 -1262
rect 1963 -1314 1973 -1262
rect 1183 -1562 1357 -1362
rect 1969 -1427 2461 -1362
rect 1969 -1484 1985 -1427
rect 2125 -1484 2461 -1427
rect 2489 -1457 2499 -1405
rect 3099 -1457 3105 -1405
rect 2489 -1473 2504 -1457
rect 3095 -1473 3105 -1457
rect 1969 -1562 2461 -1484
rect 2462 -1562 2493 -1505
rect 1353 -1662 1363 -1610
rect 1963 -1662 1973 -1610
rect 2271 -1905 2493 -1562
rect 2489 -1953 3109 -1937
rect 2489 -2005 2499 -1953
rect 3099 -2005 3109 -1953
rect 3137 -2115 3279 -718
rect 3671 -721 3793 -538
rect 3821 -673 3831 -621
rect 4431 -673 4441 -621
rect 3671 -921 3825 -721
rect 4437 -921 4591 -721
rect 3821 -1021 3831 -969
rect 4431 -1021 4438 -969
rect 4466 -1104 4591 -921
rect 3705 -1225 4591 -1104
rect 3705 -1226 4557 -1225
rect 3705 -1400 3796 -1226
rect 3824 -1352 3830 -1300
rect 4431 -1352 4441 -1300
rect 3824 -1368 4441 -1352
rect 3705 -1599 3773 -1400
rect 3825 -1599 3835 -1400
rect 3705 -1600 3824 -1599
rect 4437 -1600 4591 -1400
rect 3821 -1700 3831 -1648
rect 4432 -1700 4442 -1648
rect 3579 -1926 3589 -1848
rect 3729 -1926 3739 -1848
rect 4470 -2034 4591 -1600
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 3487 -2121 4591 -2034
rect 3487 -2244 3529 -2121
rect 4529 -2244 4591 -2121
rect 3487 -2313 4591 -2244
rect 3487 -2314 3804 -2313
<< via1 >>
rect 1363 -710 1963 -658
rect 2499 -670 3099 -618
rect 2205 -887 2345 -830
rect 1363 -1058 1963 -1006
rect 2499 -1219 3099 -1167
rect 1363 -1314 1963 -1262
rect 1985 -1484 2125 -1427
rect 2499 -1457 3099 -1405
rect 1363 -1662 1963 -1610
rect 2499 -2005 3099 -1953
rect 3831 -673 4431 -621
rect 3831 -1021 4431 -969
rect 3830 -1352 4431 -1300
rect 3773 -1599 3825 -1400
rect 3831 -1700 4432 -1648
rect 3589 -1926 3729 -1848
<< metal2 >>
rect 2499 -616 4431 -606
rect 2499 -618 3592 -616
rect 1363 -657 2135 -643
rect 1363 -658 1985 -657
rect 1963 -710 1985 -658
rect 1363 -714 1985 -710
rect 2125 -714 2135 -657
rect 3099 -670 3592 -618
rect 2499 -673 3592 -670
rect 3732 -621 4431 -616
rect 3732 -673 3831 -621
rect 2499 -683 4431 -673
rect 1363 -720 2135 -714
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -897 2355 -887
rect 3580 -969 4431 -959
rect 1363 -1006 2135 -996
rect 1963 -1058 1985 -1006
rect 1363 -1063 1985 -1058
rect 2125 -1063 2135 -1006
rect 3580 -1026 3590 -969
rect 3730 -1021 3831 -969
rect 3730 -1026 4431 -1021
rect 3580 -1036 4431 -1026
rect 1363 -1068 2135 -1063
rect 1363 -1073 2125 -1068
rect 2499 -1164 3740 -1157
rect 2499 -1167 3590 -1164
rect 3099 -1219 3590 -1167
rect 2499 -1221 3590 -1219
rect 3730 -1221 3740 -1164
rect 2499 -1229 3740 -1221
rect 1363 -1257 2355 -1247
rect 1363 -1262 2205 -1257
rect 1963 -1314 2205 -1262
rect 2345 -1314 2355 -1257
rect 1363 -1324 2355 -1314
rect 3580 -1294 4431 -1285
rect 3580 -1351 3590 -1294
rect 3730 -1300 4431 -1294
rect 3730 -1351 3830 -1300
rect 3580 -1352 3830 -1351
rect 3580 -1362 4431 -1352
rect 2499 -1400 3825 -1390
rect 2499 -1405 3177 -1400
rect 1975 -1427 2135 -1417
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 3099 -1457 3177 -1405
rect 3317 -1457 3773 -1400
rect 2499 -1467 3773 -1457
rect 1975 -1494 2135 -1484
rect 1363 -1610 2355 -1600
rect 3773 -1609 3825 -1599
rect 1963 -1662 2205 -1610
rect 1363 -1667 2205 -1662
rect 2345 -1667 2355 -1610
rect 1363 -1672 2355 -1667
rect 3580 -1648 4432 -1638
rect 3580 -1705 3590 -1648
rect 3730 -1700 3831 -1648
rect 3730 -1705 4432 -1700
rect 3580 -1715 4432 -1705
rect 3589 -1848 3729 -1838
rect 3589 -1936 3729 -1926
rect 2499 -1952 3327 -1943
rect 2499 -1953 3177 -1952
rect 3099 -2005 3177 -1953
rect 2499 -2009 3177 -2005
rect 3317 -2009 3327 -1952
rect 2499 -2015 3327 -2009
<< via2 >>
rect 1985 -714 2125 -657
rect 3592 -673 3732 -616
rect 2205 -887 2345 -830
rect 1985 -1063 2125 -1006
rect 3590 -1026 3730 -969
rect 3590 -1221 3730 -1164
rect 2205 -1314 2345 -1257
rect 3590 -1351 3730 -1294
rect 1985 -1484 2125 -1427
rect 3177 -1457 3317 -1400
rect 2205 -1667 2345 -1610
rect 3590 -1705 3730 -1648
rect 3589 -1926 3729 -1848
rect 3177 -2009 3317 -1952
<< metal3 >>
rect 3580 -616 3741 -606
rect 1975 -657 2135 -648
rect 1975 -714 1985 -657
rect 2125 -714 2135 -657
rect 1975 -1006 2135 -714
rect 3580 -673 3592 -616
rect 3732 -673 3741 -616
rect 1975 -1063 1985 -1006
rect 2125 -1063 2135 -1006
rect 1975 -1427 2135 -1063
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 1975 -1494 2135 -1484
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -1257 2355 -887
rect 2195 -1314 2205 -1257
rect 2345 -1314 2355 -1257
rect 2195 -1610 2355 -1314
rect 3580 -969 3741 -673
rect 3580 -1026 3590 -969
rect 3730 -1026 3741 -969
rect 3580 -1164 3741 -1026
rect 3580 -1221 3590 -1164
rect 3730 -1221 3741 -1164
rect 3580 -1294 3741 -1221
rect 3580 -1351 3590 -1294
rect 3730 -1351 3741 -1294
rect 2195 -1667 2205 -1610
rect 2345 -1667 2355 -1610
rect 2195 -1672 2355 -1667
rect 3167 -1400 3327 -1390
rect 3167 -1457 3177 -1400
rect 3317 -1457 3327 -1400
rect 3167 -1952 3327 -1457
rect 3580 -1648 3741 -1351
rect 3580 -1705 3590 -1648
rect 3730 -1705 3741 -1648
rect 3580 -1843 3741 -1705
rect 3579 -1848 3741 -1843
rect 3579 -1926 3589 -1848
rect 3729 -1926 3741 -1848
rect 3579 -1931 3741 -1926
rect 3167 -2009 3177 -1952
rect 3317 -2009 3327 -1952
rect 3167 -2094 3327 -2009
rect 3580 -2015 3741 -1931
use sky130_fd_pr__diode_pw2nd_05v5_37RBXE  sky130_fd_pr__diode_pw2nd_05v5_37RBXE_0
timestamp 1713020003
transform 0 1 3659 -1 0 -1887
box -183 -208 183 208
use sky130_fd_pr__nfet_01v8_MG6U6H  sky130_fd_pr__nfet_01v8_MG6U6H_0
timestamp 1713020003
transform 1 0 4131 0 1 -1500
box -496 -310 496 310
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0
timestamp 1713020003
transform -1 0 2799 0 1 -1705
box -528 -458 528 458
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1
timestamp 1713020003
transform -1 0 2799 0 1 -919
box -528 -458 528 458
use sky130_fd_pr__pfet_01v8_J2L9Q3  sky130_fd_pr__pfet_01v8_J2L9Q3_0
timestamp 1713020003
transform 1 0 4131 0 1 -821
box -496 -319 496 319
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0
timestamp 1713020003
transform 1 0 1663 0 -1 -1462
box -558 -397 558 397
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1
timestamp 1713020003
transform 1 0 1663 0 -1 -858
box -558 -397 558 397
<< labels >>
flabel space 1105 -1255 2221 -461 0 FreeSans 1600 0 0 0 M3
flabel space 2271 -1377 3327 -461 0 FreeSans 1600 0 0 0 M5
flabel space 2271 -2163 3327 -1247 0 FreeSans 1600 0 0 0 M6
flabel metal1 1183 -539 2143 -340 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 1363 -1662 1963 -1610 0 FreeSans 800 0 0 0 out_b
port 2 nsew
flabel metal2 1363 -710 1963 -658 0 FreeSans 800 0 0 0 out
port 3 nsew
flabel space 1105 -1859 2221 -1065 0 FreeSans 1600 0 0 0 M4
flabel metal1 3671 -538 4631 -340 0 FreeSans 1600 0 0 0 dvdd
port 5 nsew
flabel metal3 3580 -2015 3741 -1926 0 FreeSans 1600 0 0 0 in
port 6 nsew
flabel metal2 3317 -1467 3773 -1390 0 FreeSans 800 0 0 0 in_b
flabel metal1 2319 -2314 3279 -2115 0 FreeSans 1600 0 0 0 avss
port 4 nsew
flabel space 3635 -1810 4627 -1190 0 FreeSans 1600 0 0 0 M1
flabel space 3635 -1140 4627 -502 0 FreeSans 1600 0 0 0 M2
flabel metal1 3487 -2313 4591 -2244 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
<< end >>

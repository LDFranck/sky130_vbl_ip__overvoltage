magic
tech sky130A
magscale 1 2
timestamp 1713204736
<< metal4 >>
rect 1419 2679 1619 3382
rect 1799 2799 1999 2919
rect 1739 2739 2059 2799
rect 1679 2679 1859 2739
rect 1939 2679 2119 2739
rect 2179 2679 2379 3379
rect 1419 2619 1799 2679
rect 1999 2619 2379 2679
rect 1419 2559 1739 2619
rect 2059 2559 2379 2619
rect 1419 2499 1679 2559
rect 2119 2499 2379 2559
rect 1419 2382 1619 2499
rect 2179 2379 2379 2499
rect 2474 3179 3074 3379
rect 3195 3179 3995 3379
rect 2474 2579 2674 3179
rect 3195 2579 3395 3179
rect 3795 2579 3995 3179
rect 2474 2379 3074 2579
rect 3195 2379 3995 2579
rect 1419 1429 1619 2229
rect 2374 2029 3074 2229
rect 2474 1429 2674 2029
rect 2874 1429 3074 2029
rect 1419 1229 2019 1429
rect 2374 1229 3074 1429
rect 3395 2029 3995 2229
rect 3395 1829 3595 2029
rect 3395 1629 3895 1829
rect 3395 1229 3595 1629
rect 1419 879 2219 1079
rect 2307 879 3107 1079
rect 3195 879 3995 1079
rect 1719 79 1919 879
rect 2607 79 2807 879
rect 3495 79 3695 879
<< end >>

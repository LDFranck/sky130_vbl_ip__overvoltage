magic
tech sky130A
timestamp 1712777902
<< pwell >>
rect -164 -194 164 194
<< mvnmos >>
rect -50 -65 50 65
<< mvndiff >>
rect -79 59 -50 65
rect -79 -59 -73 59
rect -56 -59 -50 59
rect -79 -65 -50 -59
rect 50 59 79 65
rect 50 -59 56 59
rect 73 -59 79 59
rect 50 -65 79 -59
<< mvndiffc >>
rect -73 -59 -56 59
rect 56 -59 73 59
<< mvpsubdiff >>
rect -146 170 146 176
rect -146 153 -92 170
rect 92 153 146 170
rect -146 147 146 153
rect -146 122 -117 147
rect -146 -122 -140 122
rect -123 -122 -117 122
rect 117 122 146 147
rect -146 -147 -117 -122
rect 117 -122 123 122
rect 140 -122 146 122
rect 117 -147 146 -122
rect -146 -153 146 -147
rect -146 -170 -92 -153
rect 92 -170 146 -153
rect -146 -176 146 -170
<< mvpsubdiffcont >>
rect -92 153 92 170
rect -140 -122 -123 122
rect 123 -122 140 122
rect -92 -170 92 -153
<< poly >>
rect -50 101 50 109
rect -50 84 -42 101
rect 42 84 50 101
rect -50 65 50 84
rect -50 -84 50 -65
rect -50 -101 -42 -84
rect 42 -101 50 -84
rect -50 -109 50 -101
<< polycont >>
rect -42 84 42 101
rect -42 -101 42 -84
<< locali >>
rect -140 153 -92 170
rect 92 153 140 170
rect -140 122 -123 153
rect 123 122 140 153
rect -50 84 -42 101
rect 42 84 50 101
rect -73 59 -56 67
rect -73 -67 -56 -59
rect 56 59 73 67
rect 56 -67 73 -59
rect -50 -101 -42 -84
rect 42 -101 50 -84
rect -140 -153 -123 -122
rect 123 -153 140 -122
rect -140 -170 -92 -153
rect 92 -170 140 -153
<< viali >>
rect -42 84 42 101
rect -73 -59 -56 59
rect 56 -59 73 59
rect -42 -101 42 -84
<< metal1 >>
rect -48 101 48 104
rect -48 84 -42 101
rect 42 84 48 101
rect -48 81 48 84
rect -76 59 -53 65
rect -76 -59 -73 59
rect -56 -59 -53 59
rect -76 -65 -53 -59
rect 53 59 76 65
rect 53 -59 56 59
rect 73 -59 76 59
rect 53 -65 76 -59
rect -48 -84 48 -81
rect -48 -101 -42 -84
rect 42 -101 48 -84
rect -48 -104 48 -101
<< properties >>
string FIXED_BBOX -131 -161 131 161
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.3 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

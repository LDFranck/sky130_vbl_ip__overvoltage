magic
tech sky130A
magscale 1 2
timestamp 1712240559
<< pwell >>
rect -307 -1992 307 1992
<< psubdiff >>
rect -271 1922 -175 1956
rect 175 1922 271 1956
rect -271 1860 -237 1922
rect 237 1860 271 1922
rect -271 -1922 -237 -1860
rect 237 -1922 271 -1860
rect -271 -1956 -175 -1922
rect 175 -1956 271 -1922
<< psubdiffcont >>
rect -175 1922 175 1956
rect -271 -1860 -237 1860
rect 237 -1860 271 1860
rect -175 -1956 175 -1922
<< xpolycontact >>
rect -141 1394 141 1826
rect -141 -1826 141 -1394
<< xpolyres >>
rect -141 -1394 141 1394
<< locali >>
rect -271 1922 -175 1956
rect 175 1922 271 1956
rect -271 1860 -237 1922
rect 237 1860 271 1922
rect -271 -1922 -237 -1860
rect 237 -1922 271 -1860
rect -271 -1956 -175 -1922
rect 175 -1956 271 -1922
<< viali >>
rect -125 1411 125 1808
rect -125 -1808 125 -1411
<< metal1 >>
rect -131 1808 131 1820
rect -131 1411 -125 1808
rect 125 1411 131 1808
rect -131 1399 131 1411
rect -131 -1411 131 -1399
rect -131 -1808 -125 -1411
rect 125 -1808 131 -1411
rect -131 -1820 131 -1808
<< properties >>
string FIXED_BBOX -254 -1939 254 1939
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 14.1 m 1 nx 1 wmin 1.410 lmin 0.50 rho 2000 val 20.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

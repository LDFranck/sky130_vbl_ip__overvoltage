magic
tech sky130A
magscale 1 2
timestamp 1713221383
<< xpolycontact >>
rect -9024 125 -8742 557
rect -9024 -557 -8742 -125
rect -8646 125 -8364 557
rect -8646 -557 -8364 -125
rect -8268 125 -7986 557
rect -8268 -557 -7986 -125
rect -7890 125 -7608 557
rect -7890 -557 -7608 -125
rect -7512 125 -7230 557
rect -7512 -557 -7230 -125
rect -7134 125 -6852 557
rect -7134 -557 -6852 -125
rect -6756 125 -6474 557
rect -6756 -557 -6474 -125
rect -6378 125 -6096 557
rect -6378 -557 -6096 -125
rect -6000 125 -5718 557
rect -6000 -557 -5718 -125
rect -5622 125 -5340 557
rect -5622 -557 -5340 -125
rect -5244 125 -4962 557
rect -5244 -557 -4962 -125
rect -4866 125 -4584 557
rect -4866 -557 -4584 -125
rect -4488 125 -4206 557
rect -4488 -557 -4206 -125
rect -4110 125 -3828 557
rect -4110 -557 -3828 -125
rect -3732 125 -3450 557
rect -3732 -557 -3450 -125
rect -3354 125 -3072 557
rect -3354 -557 -3072 -125
rect -2976 125 -2694 557
rect -2976 -557 -2694 -125
rect -2598 125 -2316 557
rect -2598 -557 -2316 -125
rect -2220 125 -1938 557
rect -2220 -557 -1938 -125
rect -1842 125 -1560 557
rect -1842 -557 -1560 -125
rect -1464 125 -1182 557
rect -1464 -557 -1182 -125
rect -1086 125 -804 557
rect -1086 -557 -804 -125
rect -708 125 -426 557
rect -708 -557 -426 -125
rect -330 125 -48 557
rect -330 -557 -48 -125
rect 48 125 330 557
rect 48 -557 330 -125
rect 426 125 708 557
rect 426 -557 708 -125
rect 804 125 1086 557
rect 804 -557 1086 -125
rect 1182 125 1464 557
rect 1182 -557 1464 -125
rect 1560 125 1842 557
rect 1560 -557 1842 -125
rect 1938 125 2220 557
rect 1938 -557 2220 -125
rect 2316 125 2598 557
rect 2316 -557 2598 -125
rect 2694 125 2976 557
rect 2694 -557 2976 -125
rect 3072 125 3354 557
rect 3072 -557 3354 -125
rect 3450 125 3732 557
rect 3450 -557 3732 -125
rect 3828 125 4110 557
rect 3828 -557 4110 -125
rect 4206 125 4488 557
rect 4206 -557 4488 -125
rect 4584 125 4866 557
rect 4584 -557 4866 -125
rect 4962 125 5244 557
rect 4962 -557 5244 -125
rect 5340 125 5622 557
rect 5340 -557 5622 -125
rect 5718 125 6000 557
rect 5718 -557 6000 -125
rect 6096 125 6378 557
rect 6096 -557 6378 -125
rect 6474 125 6756 557
rect 6474 -557 6756 -125
rect 6852 125 7134 557
rect 6852 -557 7134 -125
rect 7230 125 7512 557
rect 7230 -557 7512 -125
rect 7608 125 7890 557
rect 7608 -557 7890 -125
rect 7986 125 8268 557
rect 7986 -557 8268 -125
rect 8364 125 8646 557
rect 8364 -557 8646 -125
rect 8742 125 9024 557
rect 8742 -557 9024 -125
<< xpolyres >>
rect -9024 -125 -8742 125
rect -8646 -125 -8364 125
rect -8268 -125 -7986 125
rect -7890 -125 -7608 125
rect -7512 -125 -7230 125
rect -7134 -125 -6852 125
rect -6756 -125 -6474 125
rect -6378 -125 -6096 125
rect -6000 -125 -5718 125
rect -5622 -125 -5340 125
rect -5244 -125 -4962 125
rect -4866 -125 -4584 125
rect -4488 -125 -4206 125
rect -4110 -125 -3828 125
rect -3732 -125 -3450 125
rect -3354 -125 -3072 125
rect -2976 -125 -2694 125
rect -2598 -125 -2316 125
rect -2220 -125 -1938 125
rect -1842 -125 -1560 125
rect -1464 -125 -1182 125
rect -1086 -125 -804 125
rect -708 -125 -426 125
rect -330 -125 -48 125
rect 48 -125 330 125
rect 426 -125 708 125
rect 804 -125 1086 125
rect 1182 -125 1464 125
rect 1560 -125 1842 125
rect 1938 -125 2220 125
rect 2316 -125 2598 125
rect 2694 -125 2976 125
rect 3072 -125 3354 125
rect 3450 -125 3732 125
rect 3828 -125 4110 125
rect 4206 -125 4488 125
rect 4584 -125 4866 125
rect 4962 -125 5244 125
rect 5340 -125 5622 125
rect 5718 -125 6000 125
rect 6096 -125 6378 125
rect 6474 -125 6756 125
rect 6852 -125 7134 125
rect 7230 -125 7512 125
rect 7608 -125 7890 125
rect 7986 -125 8268 125
rect 8364 -125 8646 125
rect 8742 -125 9024 125
<< viali >>
rect -9008 142 -8758 539
rect -8630 142 -8380 539
rect -8252 142 -8002 539
rect -7874 142 -7624 539
rect -7496 142 -7246 539
rect -7118 142 -6868 539
rect -6740 142 -6490 539
rect -6362 142 -6112 539
rect -5984 142 -5734 539
rect -5606 142 -5356 539
rect -5228 142 -4978 539
rect -4850 142 -4600 539
rect -4472 142 -4222 539
rect -4094 142 -3844 539
rect -3716 142 -3466 539
rect -3338 142 -3088 539
rect -2960 142 -2710 539
rect -2582 142 -2332 539
rect -2204 142 -1954 539
rect -1826 142 -1576 539
rect -1448 142 -1198 539
rect -1070 142 -820 539
rect -692 142 -442 539
rect -314 142 -64 539
rect 64 142 314 539
rect 442 142 692 539
rect 820 142 1070 539
rect 1198 142 1448 539
rect 1576 142 1826 539
rect 1954 142 2204 539
rect 2332 142 2582 539
rect 2710 142 2960 539
rect 3088 142 3338 539
rect 3466 142 3716 539
rect 3844 142 4094 539
rect 4222 142 4472 539
rect 4600 142 4850 539
rect 4978 142 5228 539
rect 5356 142 5606 539
rect 5734 142 5984 539
rect 6112 142 6362 539
rect 6490 142 6740 539
rect 6868 142 7118 539
rect 7246 142 7496 539
rect 7624 142 7874 539
rect 8002 142 8252 539
rect 8380 142 8630 539
rect 8758 142 9008 539
rect -9008 -539 -8758 -142
rect -8630 -539 -8380 -142
rect -8252 -539 -8002 -142
rect -7874 -539 -7624 -142
rect -7496 -539 -7246 -142
rect -7118 -539 -6868 -142
rect -6740 -539 -6490 -142
rect -6362 -539 -6112 -142
rect -5984 -539 -5734 -142
rect -5606 -539 -5356 -142
rect -5228 -539 -4978 -142
rect -4850 -539 -4600 -142
rect -4472 -539 -4222 -142
rect -4094 -539 -3844 -142
rect -3716 -539 -3466 -142
rect -3338 -539 -3088 -142
rect -2960 -539 -2710 -142
rect -2582 -539 -2332 -142
rect -2204 -539 -1954 -142
rect -1826 -539 -1576 -142
rect -1448 -539 -1198 -142
rect -1070 -539 -820 -142
rect -692 -539 -442 -142
rect -314 -539 -64 -142
rect 64 -539 314 -142
rect 442 -539 692 -142
rect 820 -539 1070 -142
rect 1198 -539 1448 -142
rect 1576 -539 1826 -142
rect 1954 -539 2204 -142
rect 2332 -539 2582 -142
rect 2710 -539 2960 -142
rect 3088 -539 3338 -142
rect 3466 -539 3716 -142
rect 3844 -539 4094 -142
rect 4222 -539 4472 -142
rect 4600 -539 4850 -142
rect 4978 -539 5228 -142
rect 5356 -539 5606 -142
rect 5734 -539 5984 -142
rect 6112 -539 6362 -142
rect 6490 -539 6740 -142
rect 6868 -539 7118 -142
rect 7246 -539 7496 -142
rect 7624 -539 7874 -142
rect 8002 -539 8252 -142
rect 8380 -539 8630 -142
rect 8758 -539 9008 -142
<< metal1 >>
rect -9014 539 -8752 551
rect -9014 142 -9008 539
rect -8758 142 -8752 539
rect -9014 130 -8752 142
rect -8636 539 -8374 551
rect -8636 142 -8630 539
rect -8380 142 -8374 539
rect -8636 130 -8374 142
rect -8258 539 -7996 551
rect -8258 142 -8252 539
rect -8002 142 -7996 539
rect -8258 130 -7996 142
rect -7880 539 -7618 551
rect -7880 142 -7874 539
rect -7624 142 -7618 539
rect -7880 130 -7618 142
rect -7502 539 -7240 551
rect -7502 142 -7496 539
rect -7246 142 -7240 539
rect -7502 130 -7240 142
rect -7124 539 -6862 551
rect -7124 142 -7118 539
rect -6868 142 -6862 539
rect -7124 130 -6862 142
rect -6746 539 -6484 551
rect -6746 142 -6740 539
rect -6490 142 -6484 539
rect -6746 130 -6484 142
rect -6368 539 -6106 551
rect -6368 142 -6362 539
rect -6112 142 -6106 539
rect -6368 130 -6106 142
rect -5990 539 -5728 551
rect -5990 142 -5984 539
rect -5734 142 -5728 539
rect -5990 130 -5728 142
rect -5612 539 -5350 551
rect -5612 142 -5606 539
rect -5356 142 -5350 539
rect -5612 130 -5350 142
rect -5234 539 -4972 551
rect -5234 142 -5228 539
rect -4978 142 -4972 539
rect -5234 130 -4972 142
rect -4856 539 -4594 551
rect -4856 142 -4850 539
rect -4600 142 -4594 539
rect -4856 130 -4594 142
rect -4478 539 -4216 551
rect -4478 142 -4472 539
rect -4222 142 -4216 539
rect -4478 130 -4216 142
rect -4100 539 -3838 551
rect -4100 142 -4094 539
rect -3844 142 -3838 539
rect -4100 130 -3838 142
rect -3722 539 -3460 551
rect -3722 142 -3716 539
rect -3466 142 -3460 539
rect -3722 130 -3460 142
rect -3344 539 -3082 551
rect -3344 142 -3338 539
rect -3088 142 -3082 539
rect -3344 130 -3082 142
rect -2966 539 -2704 551
rect -2966 142 -2960 539
rect -2710 142 -2704 539
rect -2966 130 -2704 142
rect -2588 539 -2326 551
rect -2588 142 -2582 539
rect -2332 142 -2326 539
rect -2588 130 -2326 142
rect -2210 539 -1948 551
rect -2210 142 -2204 539
rect -1954 142 -1948 539
rect -2210 130 -1948 142
rect -1832 539 -1570 551
rect -1832 142 -1826 539
rect -1576 142 -1570 539
rect -1832 130 -1570 142
rect -1454 539 -1192 551
rect -1454 142 -1448 539
rect -1198 142 -1192 539
rect -1454 130 -1192 142
rect -1076 539 -814 551
rect -1076 142 -1070 539
rect -820 142 -814 539
rect -1076 130 -814 142
rect -698 539 -436 551
rect -698 142 -692 539
rect -442 142 -436 539
rect -698 130 -436 142
rect -320 539 -58 551
rect -320 142 -314 539
rect -64 142 -58 539
rect -320 130 -58 142
rect 58 539 320 551
rect 58 142 64 539
rect 314 142 320 539
rect 58 130 320 142
rect 436 539 698 551
rect 436 142 442 539
rect 692 142 698 539
rect 436 130 698 142
rect 814 539 1076 551
rect 814 142 820 539
rect 1070 142 1076 539
rect 814 130 1076 142
rect 1192 539 1454 551
rect 1192 142 1198 539
rect 1448 142 1454 539
rect 1192 130 1454 142
rect 1570 539 1832 551
rect 1570 142 1576 539
rect 1826 142 1832 539
rect 1570 130 1832 142
rect 1948 539 2210 551
rect 1948 142 1954 539
rect 2204 142 2210 539
rect 1948 130 2210 142
rect 2326 539 2588 551
rect 2326 142 2332 539
rect 2582 142 2588 539
rect 2326 130 2588 142
rect 2704 539 2966 551
rect 2704 142 2710 539
rect 2960 142 2966 539
rect 2704 130 2966 142
rect 3082 539 3344 551
rect 3082 142 3088 539
rect 3338 142 3344 539
rect 3082 130 3344 142
rect 3460 539 3722 551
rect 3460 142 3466 539
rect 3716 142 3722 539
rect 3460 130 3722 142
rect 3838 539 4100 551
rect 3838 142 3844 539
rect 4094 142 4100 539
rect 3838 130 4100 142
rect 4216 539 4478 551
rect 4216 142 4222 539
rect 4472 142 4478 539
rect 4216 130 4478 142
rect 4594 539 4856 551
rect 4594 142 4600 539
rect 4850 142 4856 539
rect 4594 130 4856 142
rect 4972 539 5234 551
rect 4972 142 4978 539
rect 5228 142 5234 539
rect 4972 130 5234 142
rect 5350 539 5612 551
rect 5350 142 5356 539
rect 5606 142 5612 539
rect 5350 130 5612 142
rect 5728 539 5990 551
rect 5728 142 5734 539
rect 5984 142 5990 539
rect 5728 130 5990 142
rect 6106 539 6368 551
rect 6106 142 6112 539
rect 6362 142 6368 539
rect 6106 130 6368 142
rect 6484 539 6746 551
rect 6484 142 6490 539
rect 6740 142 6746 539
rect 6484 130 6746 142
rect 6862 539 7124 551
rect 6862 142 6868 539
rect 7118 142 7124 539
rect 6862 130 7124 142
rect 7240 539 7502 551
rect 7240 142 7246 539
rect 7496 142 7502 539
rect 7240 130 7502 142
rect 7618 539 7880 551
rect 7618 142 7624 539
rect 7874 142 7880 539
rect 7618 130 7880 142
rect 7996 539 8258 551
rect 7996 142 8002 539
rect 8252 142 8258 539
rect 7996 130 8258 142
rect 8374 539 8636 551
rect 8374 142 8380 539
rect 8630 142 8636 539
rect 8374 130 8636 142
rect 8752 539 9014 551
rect 8752 142 8758 539
rect 9008 142 9014 539
rect 8752 130 9014 142
rect -9014 -142 -8752 -130
rect -9014 -539 -9008 -142
rect -8758 -539 -8752 -142
rect -9014 -551 -8752 -539
rect -8636 -142 -8374 -130
rect -8636 -539 -8630 -142
rect -8380 -539 -8374 -142
rect -8636 -551 -8374 -539
rect -8258 -142 -7996 -130
rect -8258 -539 -8252 -142
rect -8002 -539 -7996 -142
rect -8258 -551 -7996 -539
rect -7880 -142 -7618 -130
rect -7880 -539 -7874 -142
rect -7624 -539 -7618 -142
rect -7880 -551 -7618 -539
rect -7502 -142 -7240 -130
rect -7502 -539 -7496 -142
rect -7246 -539 -7240 -142
rect -7502 -551 -7240 -539
rect -7124 -142 -6862 -130
rect -7124 -539 -7118 -142
rect -6868 -539 -6862 -142
rect -7124 -551 -6862 -539
rect -6746 -142 -6484 -130
rect -6746 -539 -6740 -142
rect -6490 -539 -6484 -142
rect -6746 -551 -6484 -539
rect -6368 -142 -6106 -130
rect -6368 -539 -6362 -142
rect -6112 -539 -6106 -142
rect -6368 -551 -6106 -539
rect -5990 -142 -5728 -130
rect -5990 -539 -5984 -142
rect -5734 -539 -5728 -142
rect -5990 -551 -5728 -539
rect -5612 -142 -5350 -130
rect -5612 -539 -5606 -142
rect -5356 -539 -5350 -142
rect -5612 -551 -5350 -539
rect -5234 -142 -4972 -130
rect -5234 -539 -5228 -142
rect -4978 -539 -4972 -142
rect -5234 -551 -4972 -539
rect -4856 -142 -4594 -130
rect -4856 -539 -4850 -142
rect -4600 -539 -4594 -142
rect -4856 -551 -4594 -539
rect -4478 -142 -4216 -130
rect -4478 -539 -4472 -142
rect -4222 -539 -4216 -142
rect -4478 -551 -4216 -539
rect -4100 -142 -3838 -130
rect -4100 -539 -4094 -142
rect -3844 -539 -3838 -142
rect -4100 -551 -3838 -539
rect -3722 -142 -3460 -130
rect -3722 -539 -3716 -142
rect -3466 -539 -3460 -142
rect -3722 -551 -3460 -539
rect -3344 -142 -3082 -130
rect -3344 -539 -3338 -142
rect -3088 -539 -3082 -142
rect -3344 -551 -3082 -539
rect -2966 -142 -2704 -130
rect -2966 -539 -2960 -142
rect -2710 -539 -2704 -142
rect -2966 -551 -2704 -539
rect -2588 -142 -2326 -130
rect -2588 -539 -2582 -142
rect -2332 -539 -2326 -142
rect -2588 -551 -2326 -539
rect -2210 -142 -1948 -130
rect -2210 -539 -2204 -142
rect -1954 -539 -1948 -142
rect -2210 -551 -1948 -539
rect -1832 -142 -1570 -130
rect -1832 -539 -1826 -142
rect -1576 -539 -1570 -142
rect -1832 -551 -1570 -539
rect -1454 -142 -1192 -130
rect -1454 -539 -1448 -142
rect -1198 -539 -1192 -142
rect -1454 -551 -1192 -539
rect -1076 -142 -814 -130
rect -1076 -539 -1070 -142
rect -820 -539 -814 -142
rect -1076 -551 -814 -539
rect -698 -142 -436 -130
rect -698 -539 -692 -142
rect -442 -539 -436 -142
rect -698 -551 -436 -539
rect -320 -142 -58 -130
rect -320 -539 -314 -142
rect -64 -539 -58 -142
rect -320 -551 -58 -539
rect 58 -142 320 -130
rect 58 -539 64 -142
rect 314 -539 320 -142
rect 58 -551 320 -539
rect 436 -142 698 -130
rect 436 -539 442 -142
rect 692 -539 698 -142
rect 436 -551 698 -539
rect 814 -142 1076 -130
rect 814 -539 820 -142
rect 1070 -539 1076 -142
rect 814 -551 1076 -539
rect 1192 -142 1454 -130
rect 1192 -539 1198 -142
rect 1448 -539 1454 -142
rect 1192 -551 1454 -539
rect 1570 -142 1832 -130
rect 1570 -539 1576 -142
rect 1826 -539 1832 -142
rect 1570 -551 1832 -539
rect 1948 -142 2210 -130
rect 1948 -539 1954 -142
rect 2204 -539 2210 -142
rect 1948 -551 2210 -539
rect 2326 -142 2588 -130
rect 2326 -539 2332 -142
rect 2582 -539 2588 -142
rect 2326 -551 2588 -539
rect 2704 -142 2966 -130
rect 2704 -539 2710 -142
rect 2960 -539 2966 -142
rect 2704 -551 2966 -539
rect 3082 -142 3344 -130
rect 3082 -539 3088 -142
rect 3338 -539 3344 -142
rect 3082 -551 3344 -539
rect 3460 -142 3722 -130
rect 3460 -539 3466 -142
rect 3716 -539 3722 -142
rect 3460 -551 3722 -539
rect 3838 -142 4100 -130
rect 3838 -539 3844 -142
rect 4094 -539 4100 -142
rect 3838 -551 4100 -539
rect 4216 -142 4478 -130
rect 4216 -539 4222 -142
rect 4472 -539 4478 -142
rect 4216 -551 4478 -539
rect 4594 -142 4856 -130
rect 4594 -539 4600 -142
rect 4850 -539 4856 -142
rect 4594 -551 4856 -539
rect 4972 -142 5234 -130
rect 4972 -539 4978 -142
rect 5228 -539 5234 -142
rect 4972 -551 5234 -539
rect 5350 -142 5612 -130
rect 5350 -539 5356 -142
rect 5606 -539 5612 -142
rect 5350 -551 5612 -539
rect 5728 -142 5990 -130
rect 5728 -539 5734 -142
rect 5984 -539 5990 -142
rect 5728 -551 5990 -539
rect 6106 -142 6368 -130
rect 6106 -539 6112 -142
rect 6362 -539 6368 -142
rect 6106 -551 6368 -539
rect 6484 -142 6746 -130
rect 6484 -539 6490 -142
rect 6740 -539 6746 -142
rect 6484 -551 6746 -539
rect 6862 -142 7124 -130
rect 6862 -539 6868 -142
rect 7118 -539 7124 -142
rect 6862 -551 7124 -539
rect 7240 -142 7502 -130
rect 7240 -539 7246 -142
rect 7496 -539 7502 -142
rect 7240 -551 7502 -539
rect 7618 -142 7880 -130
rect 7618 -539 7624 -142
rect 7874 -539 7880 -142
rect 7618 -551 7880 -539
rect 7996 -142 8258 -130
rect 7996 -539 8002 -142
rect 8252 -539 8258 -142
rect 7996 -551 8258 -539
rect 8374 -142 8636 -130
rect 8374 -539 8380 -142
rect 8630 -539 8636 -142
rect 8374 -551 8636 -539
rect 8752 -142 9014 -130
rect 8752 -539 8758 -142
rect 9008 -539 9014 -142
rect 8752 -551 9014 -539
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 1.41 m 1 nx 48 wmin 1.410 lmin 0.50 rho 2000 val 2.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

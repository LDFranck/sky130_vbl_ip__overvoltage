magic
tech sky130A
timestamp 1713221383
<< pwell >>
rect -264 -179 264 179
<< mvnmos >>
rect -150 -50 150 50
<< mvndiff >>
rect -179 44 -150 50
rect -179 -44 -173 44
rect -156 -44 -150 44
rect -179 -50 -150 -44
rect 150 44 179 50
rect 150 -44 156 44
rect 173 -44 179 44
rect 150 -50 179 -44
<< mvndiffc >>
rect -173 -44 -156 44
rect 156 -44 173 44
<< mvpsubdiff >>
rect -246 155 246 161
rect -246 138 -192 155
rect 192 138 246 155
rect -246 132 246 138
rect -246 107 -217 132
rect -246 -107 -240 107
rect -223 -107 -217 107
rect 217 107 246 132
rect -246 -132 -217 -107
rect 217 -107 223 107
rect 240 -107 246 107
rect 217 -132 246 -107
rect -246 -138 246 -132
rect -246 -155 -192 -138
rect 192 -155 246 -138
rect -246 -161 246 -155
<< mvpsubdiffcont >>
rect -192 138 192 155
rect -240 -107 -223 107
rect 223 -107 240 107
rect -192 -155 192 -138
<< poly >>
rect -150 86 150 94
rect -150 69 -142 86
rect 142 69 150 86
rect -150 50 150 69
rect -150 -69 150 -50
rect -150 -86 -142 -69
rect 142 -86 150 -69
rect -150 -94 150 -86
<< polycont >>
rect -142 69 142 86
rect -142 -86 142 -69
<< locali >>
rect -240 138 -192 155
rect 192 138 240 155
rect -240 107 -223 138
rect 223 107 240 138
rect -150 69 -142 86
rect 142 69 150 86
rect -173 44 -156 52
rect -173 -52 -156 -44
rect 156 44 173 52
rect 156 -52 173 -44
rect -150 -86 -142 -69
rect 142 -86 150 -69
rect -240 -138 -223 -107
rect 223 -138 240 -107
rect -240 -155 -192 -138
rect 192 -155 240 -138
<< viali >>
rect -142 69 142 86
rect -173 -44 -156 44
rect 156 -44 173 44
rect -142 -86 142 -69
<< metal1 >>
rect -148 86 148 89
rect -148 69 -142 86
rect 142 69 148 86
rect -148 66 148 69
rect -176 44 -153 50
rect -176 -44 -173 44
rect -156 -44 -153 44
rect -176 -50 -153 -44
rect 153 44 176 50
rect 153 -44 156 44
rect 173 -44 176 44
rect 153 -50 176 -44
rect -148 -69 148 -66
rect -148 -86 -142 -69
rect 142 -86 148 -69
rect -148 -89 148 -86
<< properties >>
string FIXED_BBOX -231 -146 231 146
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 3 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
timestamp 1712777902
<< pwell >>
rect -148 -255 148 255
<< nmos >>
rect -50 -150 50 150
<< ndiff >>
rect -79 144 -50 150
rect -79 -144 -73 144
rect -56 -144 -50 144
rect -79 -150 -50 -144
rect 50 144 79 150
rect 50 -144 56 144
rect 73 -144 79 144
rect 50 -150 79 -144
<< ndiffc >>
rect -73 -144 -56 144
rect 56 -144 73 144
<< psubdiff >>
rect -130 220 -82 237
rect 82 220 130 237
rect -130 189 -113 220
rect 113 189 130 220
rect -130 -220 -113 -189
rect 113 -220 130 -189
rect -130 -237 -82 -220
rect 82 -237 130 -220
<< psubdiffcont >>
rect -82 220 82 237
rect -130 -189 -113 189
rect 113 -189 130 189
rect -82 -237 82 -220
<< poly >>
rect -50 186 50 194
rect -50 169 -42 186
rect 42 169 50 186
rect -50 150 50 169
rect -50 -169 50 -150
rect -50 -186 -42 -169
rect 42 -186 50 -169
rect -50 -194 50 -186
<< polycont >>
rect -42 169 42 186
rect -42 -186 42 -169
<< locali >>
rect -130 220 -82 237
rect 82 220 130 237
rect -130 189 -113 220
rect 113 189 130 220
rect -50 169 -42 186
rect 42 169 50 186
rect -73 144 -56 152
rect -73 -152 -56 -144
rect 56 144 73 152
rect 56 -152 73 -144
rect -50 -186 -42 -169
rect 42 -186 50 -169
rect -130 -220 -113 -189
rect 113 -220 130 -189
rect -130 -237 -82 -220
rect 82 -237 130 -220
<< viali >>
rect -42 169 42 186
rect -73 -144 -56 144
rect 56 -144 73 144
rect -42 -186 42 -169
<< metal1 >>
rect -48 186 48 189
rect -48 169 -42 186
rect 42 169 48 186
rect -48 166 48 169
rect -76 144 -53 150
rect -76 -144 -73 144
rect -56 -144 -53 144
rect -76 -150 -53 -144
rect 53 144 76 150
rect 53 -144 56 144
rect 73 -144 76 144
rect 53 -150 76 -144
rect -48 -169 48 -166
rect -48 -186 -42 -169
rect 42 -186 48 -169
rect -48 -189 48 -186
<< properties >>
string FIXED_BBOX -121 -228 121 228
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 3.0 l 1.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

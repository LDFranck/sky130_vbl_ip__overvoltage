magic
tech sky130A
magscale 1 2
timestamp 1712073957
<< nwell >>
rect -3425 -319 3425 319
<< pmos >>
rect -3229 -100 -29 100
rect 29 -100 3229 100
<< pdiff >>
rect -3287 88 -3229 100
rect -3287 -88 -3275 88
rect -3241 -88 -3229 88
rect -3287 -100 -3229 -88
rect -29 88 29 100
rect -29 -88 -17 88
rect 17 -88 29 88
rect -29 -100 29 -88
rect 3229 88 3287 100
rect 3229 -88 3241 88
rect 3275 -88 3287 88
rect 3229 -100 3287 -88
<< pdiffc >>
rect -3275 -88 -3241 88
rect -17 -88 17 88
rect 3241 -88 3275 88
<< nsubdiff >>
rect -3389 249 -3293 283
rect 3293 249 3389 283
rect -3389 187 -3355 249
rect 3355 187 3389 249
rect -3389 -249 -3355 -187
rect 3355 -249 3389 -187
rect -3389 -283 -3293 -249
rect 3293 -283 3389 -249
<< nsubdiffcont >>
rect -3293 249 3293 283
rect -3389 -187 -3355 187
rect 3355 -187 3389 187
rect -3293 -283 3293 -249
<< poly >>
rect -3229 181 -29 197
rect -3229 147 -3213 181
rect -45 147 -29 181
rect -3229 100 -29 147
rect 29 181 3229 197
rect 29 147 45 181
rect 3213 147 3229 181
rect 29 100 3229 147
rect -3229 -147 -29 -100
rect -3229 -181 -3213 -147
rect -45 -181 -29 -147
rect -3229 -197 -29 -181
rect 29 -147 3229 -100
rect 29 -181 45 -147
rect 3213 -181 3229 -147
rect 29 -197 3229 -181
<< polycont >>
rect -3213 147 -45 181
rect 45 147 3213 181
rect -3213 -181 -45 -147
rect 45 -181 3213 -147
<< locali >>
rect -3389 249 -3293 283
rect 3293 249 3389 283
rect -3389 187 -3355 249
rect 3355 187 3389 249
rect -3229 147 -3213 181
rect -45 147 -29 181
rect 29 147 45 181
rect 3213 147 3229 181
rect -3275 88 -3241 104
rect -3275 -104 -3241 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 3241 88 3275 104
rect 3241 -104 3275 -88
rect -3229 -181 -3213 -147
rect -45 -181 -29 -147
rect 29 -181 45 -147
rect 3213 -181 3229 -147
rect -3389 -249 -3355 -187
rect 3355 -249 3389 -187
rect -3389 -283 -3293 -249
rect 3293 -283 3389 -249
<< viali >>
rect -3213 147 -45 181
rect 45 147 3213 181
rect -3275 -88 -3241 88
rect -17 -88 17 88
rect 3241 -88 3275 88
rect -3213 -181 -45 -147
rect 45 -181 3213 -147
<< metal1 >>
rect -3225 181 -33 187
rect -3225 147 -3213 181
rect -45 147 -33 181
rect -3225 141 -33 147
rect 33 181 3225 187
rect 33 147 45 181
rect 3213 147 3225 181
rect 33 141 3225 147
rect -3281 88 -3235 100
rect -3281 -88 -3275 88
rect -3241 -88 -3235 88
rect -3281 -100 -3235 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 3235 88 3281 100
rect 3235 -88 3241 88
rect 3275 -88 3281 88
rect 3235 -100 3281 -88
rect -3225 -147 -33 -141
rect -3225 -181 -3213 -147
rect -45 -181 -33 -147
rect -3225 -187 -33 -181
rect 33 -147 3225 -141
rect 33 -181 45 -147
rect 3213 -181 3225 -147
rect 33 -187 3225 -181
<< properties >>
string FIXED_BBOX -3372 -266 3372 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 16 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

* PEX produced on dom 21 abr 2024 23:23:20 -03 using ./iic-pex.sh with m=3 and s=1
* NGSPICE file created from sky130_vbl_ip__overvoltage.ext - technology: sky130A

.subckt sky130_vbl_ip__overvoltage vtrip[3] vtrip[2] ovout vtrip[0] vbg ibias ena
+ vtrip[1] dvss dvdd avdd avss
X0 dvss.t73 dvss.t71 dvss.t72 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X1 multiplexer_0.trans_gate_m_31.out.t4 multiplexer_0.vtrip_1.t2 multiplexer_0.trans_gate_m_29.in.t5 avss.t217 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X2 avss.t44 multiplexer_0.vtrip_1_b.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X3 a_n15874_n447.t1 a_n12654_n447.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X4 a_n12118_12027.t1 a_n8898_11649.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X5 dvss.t70 dvss.t68 dvss.t69 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X6 avss.t218 avss.t219 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X7 avss.t33 avss.t34 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X8 comp_hyst_0.net3.t3 comp_hyst_0.net4.t11 dvdd.t12 dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X9 avss.t19 avss.t20 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X10 avss.t88 avss.t89 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X11 avss.t247 level_shifter_3.in_b.t2 multiplexer_0.vtrip_3.t1 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X12 a_n8362_4845.t0 multiplexer_0.in_0110.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X13 a_n15874_8625.t1 a_n12654_9003.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X14 avss.t131 multiplexer_0.vtrip_2.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X15 a_n12118_9759.t0 a_n8898_9381.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X16 multiplexer_0.in_1100.t0 multiplexer_0.in_1101.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X17 dvss.t67 dvss.t65 dvss.t66 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X18 a_n15874_6357.t0 a_n12654_5979.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X19 level_shifter_0.in_b.t0 vtrip[0].t0 dvdd.t5 dvdd.t4 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X20 dvdd.t113 dvdd.t111 dvdd.t112 dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X21 multiplexer_0.trans_gate_m_37.out.t5 multiplexer_0.vtrip_2.t3 multiplexer_0.trans_gate_m_32.in.t3 avdd.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X22 multiplexer_0.trans_gate_m_21.in.t0 multiplexer_0.vtrip_0.t2 multiplexer_0.in_1011.t0 avss.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X23 avss.t142 vtrip[1].t0 multiplexer_0.vtrip_1_b.t0 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X24 dvss.t20 comp_hyst_0.net5.t5 comp_hyst_0.net1.t0 dvss.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X25 avss.t172 avss.t173 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X26 multiplexer_0.trans_gate_m_29.in.t1 multiplexer_0.vtrip_0.t3 multiplexer_0.in_0010.t0 avdd.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X27 avss.t73 multiplexer_0.vtrip_0_b.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X28 a_n12118_2955.t1 a_n8898_3333.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X29 avss.t212 avss.t213 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X30 avss.t127 avss.t128 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X31 voltage_divider_0.51.t1 multiplexer_0.in_0000.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X32 avss.t42 avss.t43 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X33 comp_hyst_0.net1.t1 vin.t4 comp_hyst_0.net3.t0 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X34 a_n15874_13161.t0 a_n12654_13539.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X35 multiplexer_0.trans_gate_m_23.in.t3 multiplexer_0.vtrip_0_b.t3 multiplexer_0.in_1001.t3 avdd.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X36 a_n8362_13161.t0 a_n5142_12783.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X37 avss.t170 avss.t171 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X38 avss.t95 avss.t96 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X39 a_n12118_7491.t0 a_n8898_7113.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X40 multiplexer_0.trans_gate_m_32.in.t1 multiplexer_0.vtrip_1.t3 multiplexer_0.trans_gate_m_23.in.t2 avdd.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X41 multiplexer_0.vtrip_2.t0 multiplexer_0.vtrip_2_b.t2 avdd.t2 avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X42 avss.t99 avss.t100 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X43 dvdd.t110 dvdd.t108 dvdd.t109 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X44 a_n15874_3333.t0 a_n12654_3711.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X45 a_n8898_n447.t1 a_n5142_n825.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X46 comp_hyst_0.net1.t3 vbg.t0 comp_hyst_0.net4.t8 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X47 avss.t168 avss.t169 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X48 avss.t84 avss.t85 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X49 avss.t185 level_shifter_0.in_b.t2 multiplexer_0.vtrip_0.t1 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X50 a_n12118_10515.t1 a_n8898_10893.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X51 comp_hyst_0.net4.t10 comp_hyst_0.net3.t9 dvdd.t120 dvdd.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X52 a_n8362_8625.t0 multiplexer_0.in_0000.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X53 multiplexer_0.in_0100.t0 a_n5142_5979.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X54 dvdd.t107 dvdd.t105 dvdd.t106 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X55 a_n15874_10893.t1 a_n12654_11271.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X56 comp_hyst_0.net1.t2 vin.t5 comp_hyst_0.net3.t1 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X57 multiplexer_0.trans_gate_m_27.in.t1 multiplexer_0.vtrip_0.t4 multiplexer_0.in_0101.t0 avss.t191 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X58 avss.t74 avss.t75 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X59 comp_hyst_0.net1.t4 vbg.t1 comp_hyst_0.net4.t9 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
X60 avss.t125 avss.t126 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X61 a_n8362_10137.t1 a_n5142_9759.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X62 a_n12118_6735.t0 a_n8898_7113.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X63 multiplexer_0.trans_gate_m_28.in.t5 multiplexer_0.vtrip_1_b.t3 multiplexer_0.trans_gate_m_27.in.t5 avss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X64 avss.t81 ena.t0 a_n5142_n1959.t0 avss.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=3
X65 dvdd.t104 dvdd.t102 dvdd.t103 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X66 a_n12118_4467.t1 a_n8898_4089.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X67 avss.t82 avss.t83 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X68 dvss.t64 dvss.t62 dvss.t63 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X69 a_n15874_1065.t0 a_n12654_1065.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X70 multiplexer_0.vtrip_3.t0 multiplexer_0.vtrip_3_b.t2 avdd.t27 avdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X71 vin.t3 multiplexer_0.vtrip_3_b.t3 multiplexer_0.trans_gate_m_33.in.t2 avss.t246 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X72 avss.t189 multiplexer_0.vtrip_1_b.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X73 avss.t123 avss.t124 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X74 a_n8362_13917.t0 a_n5142_14295.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X75 dvdd.t101 dvdd.t99 dvdd.t100 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X76 multiplexer_0.trans_gate_m_33.in.t5 multiplexer_0.vtrip_2.t4 multiplexer_0.trans_gate_m_31.out.t5 avdd.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X77 avss.t208 avss.t209 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X78 a_n12118_10515.t0 a_n8898_10137.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X79 avss.t202 avss.t203 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X80 a_n8362_13917.t1 a_n5142_13539.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X81 multiplexer_0.in_1010.t1 multiplexer_0.in_1001.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X82 a_n15874_n447.t0 a_n12654_n69.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X83 a_n15874_4845.t1 a_n12654_4467.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X84 avss.t121 avss.t122 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X85 dvss.t24 comp_hyst_0.ena_b.t2 comp_hyst_0.net5.t3 dvss.t23 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X86 a_n12118_14295.t0 a_n8898_14673.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X87 level_shifter_2.in_b.t0 vtrip[2].t0 dvdd.t117 dvdd.t116 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X88 dvdd.t98 dvdd.t96 dvdd.t97 dvdd.t53 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X89 a_n12654_1821.t1 a_n8898_1821.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X90 a_n15874_14673.t0 a_n12654_15051.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X91 avss.t210 avss.t211 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X92 multiplexer_0.trans_gate_m_18.in.t1 multiplexer_0.vtrip_0.t5 multiplexer_0.in_1100.t3 avdd.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X93 avss.t54 level_shifter_2.in_b.t2 multiplexer_0.vtrip_2.t1 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X94 avss.t93 avss.t94 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X95 multiplexer_0.trans_gate_m_32.in.t4 multiplexer_0.vtrip_1_b.t5 multiplexer_0.trans_gate_m_21.in.t5 avdd.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X96 comp_hyst_0.net3.t7 comp_hyst_0.net3.t6 dvdd.t20 dvdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X97 avss.t119 avss.t120 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X98 dvss.t22 vtrip[2].t1 level_shifter_2.in_b.t1 dvss.t21 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X99 a_n12118_8247.t0 a_n8898_7869.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X100 multiplexer_0.trans_gate_m_19.in.t3 multiplexer_0.vtrip_0_b.t4 multiplexer_0.in_1110.t3 avss.t197 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X101 dvss.t16 comp_hyst_0.net2 comp_hyst_0.net2.t2 dvss.t15 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X102 a_n15874_n1959.t0 a_n12654_n1959.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X103 a_n8898_1065.t0 a_n5142_687.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X104 multiplexer_0.vtrip_0_b.t0 multiplexer_0.vtrip_0.t6 avdd.t14 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X105 multiplexer_0.trans_gate_m_29.in.t4 multiplexer_0.vtrip_0_b.t5 multiplexer_0.in_0011.t3 avdd.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X106 avss.t71 avss.t72 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X107 multiplexer_0.trans_gate_m_33.in.t4 multiplexer_0.vtrip_2.t5 multiplexer_0.trans_gate_m_28.in.t3 avss.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X108 avss.t44 multiplexer_0.vtrip_1.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X109 dvdd.t95 dvdd.t93 dvdd.t94 dvdd.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X110 a_n8898_n1581.t1 a_n5142_n1581.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X111 a_n15874_1821.t1 a_n12654_2199.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X112 a_n12654_n69.t0 a_n8898_n69.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X113 a_n12118_11271.t0 a_n8898_11649.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X114 avss.t183 avss.t184 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X115 a_n8362_4845.t1 multiplexer_0.in_0111.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X116 a_n15874_11649.t1 a_n12654_12027.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X117 a_n15874_8625.t0 a_n12654_8247.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X118 avss.t255 avss.t256 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X119 multiplexer_0.trans_gate_m_19.in.t1 multiplexer_0.vtrip_0.t7 multiplexer_0.in_1111.t0 avss.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X120 avss.t200 avss.t201 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X121 a_n15874_5601.t0 a_n12654_5979.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X122 avss.t73 multiplexer_0.vtrip_0.t8 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X123 multiplexer_0.trans_gate_m_28.in.t1 multiplexer_0.vtrip_1.t5 multiplexer_0.trans_gate_m_25.in.t2 avss.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X124 comp_hyst_0.net4.t5 comp_hyst_0.net3.t10 dvdd.t17 dvdd.t16 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X125 avss.t52 avss.t53 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X126 avss.t69 avss.t70 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X127 multiplexer_0.trans_gate_m_37.in.t2 multiplexer_0.vtrip_1.t6 multiplexer_0.trans_gate_m_19.in.t2 avss.t215 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X128 a_n12118_5223.t1 a_n8898_5601.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X129 a_n8898_n1203.t1 a_n5142_n1581.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X130 a_n12118_2955.t0 a_n8898_2577.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X131 avss.t110 avss.t111 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X132 multiplexer_0.trans_gate_m_25.in.t3 multiplexer_0.vtrip_0_b.t6 multiplexer_0.in_0111.t3 avdd.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X133 dvdd.t92 dvdd.t90 dvdd.t91 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X134 avss.t117 avss.t118 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X135 comp_hyst_0.net4.t0 ena.t1 dvdd.t3 dvdd.t2 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X136 avss.t11 avss.t12 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X137 a_n8362_12405.t0 a_n5142_12783.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X138 multiplexer_0.trans_gate_m_23.in.t4 multiplexer_0.vtrip_0_b.t7 multiplexer_0.in_1000.t3 avss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X139 multiplexer_0.trans_gate_m_37.out.t1 multiplexer_0.vtrip_2_b.t3 multiplexer_0.trans_gate_m_37.in.t0 avdd.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X140 avss.t152 ena.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X141 dvdd.t89 dvdd.t87 dvdd.t88 dvdd.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X142 multiplexer_0.in_1110.t2 multiplexer_0.in_1101.t3 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X143 dvdd.t86 dvdd.t84 dvdd.t85 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X144 multiplexer_0.vtrip_3_b.t0 multiplexer_0.vtrip_3.t2 avdd.t25 avdd.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X145 comp_hyst_0.net2.t0 comp_hyst_0.net4.t12 dvdd.t11 dvdd.t10 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X146 vin.t2 multiplexer_0.vtrip_3.t3 multiplexer_0.trans_gate_m_37.out.t3 avss.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X147 avss.t166 avss.t167 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X148 multiplexer_0.trans_gate_m_27.in.t0 multiplexer_0.vtrip_0.t9 multiplexer_0.in_0100.t1 avdd.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X149 avss.t91 avss.t92 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X150 avss.t58 avss.t59 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X151 avss.t250 avss.t251 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X152 multiplexer_0.trans_gate_m_31.in.t1 multiplexer_0.vtrip_0.t10 multiplexer_0.in_0000.t0 avdd.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X153 a_n8362_8625.t1 multiplexer_0.in_0001.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X154 avss.t67 avss.t68 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X155 multiplexer_0.in_0101.t2 a_n5142_5979.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X156 multiplexer_0.trans_gate_m_37.in.t1 multiplexer_0.vtrip_1.t7 multiplexer_0.trans_gate_m_18.in.t2 avdd.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X157 a_n12654_n825.t1 a_n8898_n825.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X158 avss.t232 avss.t233 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X159 a_n15874_9381.t0 a_n12654_9759.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X160 a_n15874_10893.t0 a_n12654_10515.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X161 avss.t198 avss.t199 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X162 a_n8362_12405.t1 a_n5142_12027.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X163 dvss.t18 vbg.t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X164 a_n12118_6735.t1 a_n8898_6357.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X165 avss.t164 avss.t165 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X166 a_n15874_3333.t1 a_n12654_2955.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X167 avss.t27 avss.t28 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X168 avss.t248 avss.t249 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X169 a_n12118_12783.t1 a_n8898_13161.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X170 multiplexer_0.trans_gate_m_18.in.t3 multiplexer_0.vtrip_0_b.t8 multiplexer_0.in_1101.t0 avdd.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X171 dvss.t26 comp_hyst_0.ena_b.t3 comp_hyst_0.net2.t1 dvss.t25 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X172 dvdd.t83 dvdd.t81 dvdd.t82 dvdd.t53 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X173 multiplexer_0.trans_gate_m_31.out.t3 multiplexer_0.vtrip_1.t8 multiplexer_0.trans_gate_m_31.in.t2 avdd.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X174 a_n15874_7113.t1 a_n12654_7491.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X175 comp_hyst_0.ena_b.t0 ena.t3 dvdd.t115 dvdd.t114 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X176 a_n15874_10137.t1 a_n12654_10515.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X177 avss.t55 avss.t56 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X178 multiplexer_0.trans_gate_m_37.out.t0 multiplexer_0.vtrip_2_b.t4 multiplexer_0.trans_gate_m_32.in.t0 avss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X179 multiplexer_0.vtrip_1.t1 multiplexer_0.vtrip_1_b.t6 avdd.t39 avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X180 avss.t194 avss.t195 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X181 multiplexer_0.trans_gate_m_29.in.t0 multiplexer_0.vtrip_0_b.t9 multiplexer_0.in_0010.t2 avss.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X182 dvdd.t80 dvdd.t78 dvdd.t79 dvdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X183 a_n12118_3711.t0 a_n8898_4089.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X184 avss.t161 multiplexer_0.vtrip_3_b.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X185 avss.t230 avss.t231 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X186 avss.t149 avss.t150 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X187 avss.t238 vtrip[3].t0 multiplexer_0.vtrip_3_b.t1 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X188 a_n15874_309.t0 a_n12654_687.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X189 voltage_divider_0.51.t0 a_n5142_9759.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X190 a_n15874_14673.t1 a_n12654_14295.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X191 dvdd.t77 dvdd.t75 dvdd.t76 dvdd.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X192 dvss.t28 ena.t4 comp_hyst_0.ena_b.t1 dvss.t27 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X193 multiplexer_0.trans_gate_m_23.in.t0 multiplexer_0.vtrip_0.t11 multiplexer_0.in_1001.t0 avss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X194 comp_hyst_0.net5.t4 ena.t5 ibias.t0 dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
X195 a_n12118_9759.t1 a_n8898_10137.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X196 avss.t244 avss.t245 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X197 a_n8362_13161.t1 a_n5142_13539.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X198 multiplexer_0.trans_gate_m_32.in.t5 multiplexer_0.vtrip_1_b.t7 multiplexer_0.trans_gate_m_23.in.t5 avss.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X199 multiplexer_0.in_1010.t2 multiplexer_0.in_1011.t3 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X200 a_n15874_7113.t0 a_n12654_6735.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X201 a_n12118_7491.t1 a_n8898_7869.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X202 a_n15874_4089.t0 a_n12654_4467.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X203 avss.t45 avss.t46 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X204 dvss.t74 ena.t6 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X205 a_n12118_14295.t1 a_n8898_13917.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X206 level_shifter_1.in_b.t0 vtrip[1].t1 dvdd.t22 dvdd.t21 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X207 dvdd.t74 dvdd.t72 dvdd.t73 dvdd.t16 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X208 avss.t6 avss.t7 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X209 multiplexer_0.trans_gate_m_21.in.t1 multiplexer_0.vtrip_0.t12 multiplexer_0.in_1010.t0 avdd.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X210 dvdd.t71 dvdd.t69 dvdd.t70 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X211 multiplexer_0.trans_gate_m_28.in.t2 multiplexer_0.vtrip_1.t9 multiplexer_0.trans_gate_m_27.in.t2 avdd.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X212 a_n12118_13539.t1 a_n8898_13917.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X213 a_n12654_1443.t0 a_n8898_1443.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X214 a_n8362_7113.t1 multiplexer_0.in_0010.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X215 avss.t192 avss.t193 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X216 avss.t32 level_shifter_1.in_b.t2 multiplexer_0.vtrip_1.t0 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X217 a_n15874_309.t1 a_n12654_309.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X218 a_n8898_n69.t1 a_n5142_n69.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X219 avss.t17 avss.t18 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X220 a_n12654_687.t0 a_n8898_687.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X221 a_n15874_11649.t0 a_n12654_11271.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X222 dvdd.t68 dvdd.t66 dvdd.t67 dvdd.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X223 dvss.t12 vtrip[3].t1 level_shifter_3.in_b.t1 dvss.t11 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X224 dvdd.t65 dvdd.t63 dvdd.t64 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X225 a_n8362_10893.t0 a_n5142_11271.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X226 avss.t242 avss.t243 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X227 avss.t139 avss.t140 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X228 multiplexer_0.trans_gate_m_18.in.t0 multiplexer_0.vtrip_0.t13 multiplexer_0.in_1101.t1 avss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X229 avss.t155 avss.t156 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X230 dvss.t7 vtrip[1].t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X231 avss.t115 avss.t116 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X232 dvdd.t62 dvdd.t59 dvdd.t61 dvdd.t60 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X233 a_n15874_1821.t0 a_n12654_1821.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X234 comp_hyst_0.net4.t6 comp_hyst_0.net3.t11 dvdd.t19 dvdd.t18 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X235 multiplexer_0.trans_gate_m_31.in.t4 multiplexer_0.vtrip_0_b.t10 multiplexer_0.in_0001.t3 avdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X236 avss.t162 avss.t163 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X237 multiplexer_0.trans_gate_m_25.in.t4 multiplexer_0.vtrip_0_b.t11 multiplexer_0.in_0110.t2 avss.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X238 avss.t240 avss.t241 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X239 multiplexer_0.trans_gate_m_33.in.t1 multiplexer_0.vtrip_2_b.t5 multiplexer_0.trans_gate_m_31.out.t0 avss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X240 multiplexer_0.trans_gate_m_37.in.t5 multiplexer_0.vtrip_1_b.t8 multiplexer_0.trans_gate_m_19.in.t5 avdd.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X241 avss.t236 avss.t237 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X242 a_n8362_7113.t0 multiplexer_0.in_0011.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X243 a_n12654_n1581.t1 a_n8898_n1581.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X244 multiplexer_0.in_1000.t2 multiplexer_0.in_0111.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X245 a_n15874_7869.t1 a_n12654_8247.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X246 dvss.t9 vtrip[1].t3 level_shifter_1.in_b.t1 dvss.t8 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X247 a_n12654_309.t0 a_n8898_309.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X248 comp_hyst_0.net4.t2 comp_hyst_0.net4.t1 dvdd.t9 dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X249 avss.t90 vtrip[0].t1 multiplexer_0.vtrip_0_b.t1 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X250 avss.t50 avss.t51 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X251 avss.t48 avss.t49 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X252 a_n12118_5223.t0 a_n8898_4845.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X253 a_n12118_2199.t1 a_n8898_2577.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X254 level_shifter_3.in_b.t0 vtrip[3].t2 dvdd.t1 dvdd.t0 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X255 avss.t180 avss.t181 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X256 dvdd.t58 dvdd.t56 dvdd.t57 dvdd.t53 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X257 multiplexer_0.trans_gate_m_31.out.t1 multiplexer_0.vtrip_1_b.t9 multiplexer_0.trans_gate_m_29.in.t3 avdd.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X258 avss.t147 multiplexer_0.vtrip_0.t14 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X259 a_n8898_15051.t1 avdd.t28 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X260 avss.t234 avss.t235 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X261 avss.t23 avss.t24 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X262 avss.t137 avss.t138 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X263 avss.t178 avss.t179 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X264 multiplexer_0.trans_gate_m_32.in.t2 multiplexer_0.vtrip_1.t10 multiplexer_0.trans_gate_m_21.in.t3 avss.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X265 avss.t176 avss.t177 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X266 a_n12118_9003.t1 a_n8898_9381.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X267 avss.t3 avss.t4 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X268 a_n12654_n1203.t1 a_n8898_n1203.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X269 multiplexer_0.trans_gate_m_29.in.t2 multiplexer_0.vtrip_0.t15 multiplexer_0.in_0011.t0 avss.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X270 dvdd.t55 dvdd.t52 dvdd.t54 dvdd.t53 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X271 multiplexer_0.in_1110.t1 multiplexer_0.in_1111.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X272 dvdd.t51 dvdd.t49 dvdd.t50 dvdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X273 a_n15874_5601.t1 a_n12654_5223.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X274 multiplexer_0.vtrip_2_b.t1 multiplexer_0.vtrip_2.t6 avdd.t29 avdd.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X275 a_n15874_2577.t0 a_n12654_2955.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X276 multiplexer_0.trans_gate_m_21.in.t2 multiplexer_0.vtrip_0_b.t12 multiplexer_0.in_1011.t2 avdd.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X277 a_n8898_n1959.t1 a_n5142_n1959.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X278 dvdd.t48 dvdd.t46 dvdd.t47 dvdd.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X279 avss.t113 avss.t114 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X280 a_n12118_12783.t0 a_n8898_12405.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X281 multiplexer_0.trans_gate_m_18.in.t4 multiplexer_0.vtrip_0_b.t13 multiplexer_0.in_1100.t2 avss.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X282 dvss.t17 vtrip[3].t3 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X283 a_n8362_7869.t1 multiplexer_0.in_0001.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X284 a_n15874_13161.t1 a_n12654_12783.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X285 comp_hyst_0.net3.t5 comp_hyst_0.net3.t4 dvdd.t14 dvdd.t13 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X286 ovout.t2 comp_hyst_0.net3.t12 dvdd.t24 dvdd.t23 sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
X287 a_n12654_n447.t0 a_n8898_n447.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X288 avss.t108 avss.t109 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X289 dvdd.t45 dvdd.t42 dvdd.t44 dvdd.t43 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X290 a_n8362_11649.t0 a_n5142_12027.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X291 avss.t190 multiplexer_0.vtrip_3.t4 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X292 avss.t97 avss.t98 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X293 a_n12118_9003.t0 a_n8898_8625.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X294 a_n12118_5979.t0 a_n8898_6357.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X295 dvdd.t41 dvdd.t39 dvdd.t40 dvdd.t16 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=16
X296 avss.t106 avss.t107 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X297 multiplexer_0.trans_gate_m_25.in.t0 multiplexer_0.vtrip_0.t16 multiplexer_0.in_0111.t0 avss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X298 dvdd.t38 dvdd.t36 dvdd.t37 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X299 a_n15874_n1203.t0 a_n12654_n825.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X300 avss.t15 avss.t16 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X301 a_n12118_12027.t0 a_n8898_12405.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X302 avss.t1 avss.t2 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X303 comp_hyst_0.net4.t7 comp_hyst_0.net3.t13 dvdd.t25 dvdd.t16 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
X304 avss.t21 avss.t22 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X305 multiplexer_0.in_0101.t1 multiplexer_0.in_0110.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X306 avss.t104 avss.t105 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X307 a_n15874_10137.t0 a_n12654_9759.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X308 multiplexer_0.vtrip_0.t0 multiplexer_0.vtrip_0_b.t14 avdd.t32 avdd.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X309 multiplexer_0.in_1100.t1 multiplexer_0.in_1011.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X310 a_n15874_6357.t1 a_n12654_6735.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X311 multiplexer_0.trans_gate_m_27.in.t4 multiplexer_0.vtrip_0_b.t15 multiplexer_0.in_0101.t3 avdd.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X312 avss.t226 avss.t227 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X313 avss.t66 vtrip[2].t2 multiplexer_0.vtrip_2_b.t0 avss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
X314 a_n12118_3711.t1 a_n8898_3333.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X315 dvss.t61 dvss.t59 dvss.t60 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X316 multiplexer_0.trans_gate_m_31.in.t3 multiplexer_0.vtrip_0_b.t16 multiplexer_0.in_0000.t3 avss.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X317 avss.t206 avss.t207 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X318 a_n15874_13917.t1 a_n12654_14295.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X319 vin.t1 multiplexer_0.vtrip_3.t5 multiplexer_0.trans_gate_m_33.in.t3 avdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X320 avss.t224 avss.t225 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X321 a_n15874_13917.t0 a_n12654_13539.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X322 avss.t222 avss.t223 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X323 avss.t220 avss.t221 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X324 multiplexer_0.trans_gate_m_37.out.t4 multiplexer_0.vtrip_2.t7 multiplexer_0.trans_gate_m_37.in.t3 avss.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X325 dvss.t6 vin.t6 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X326 a_n8362_10893.t1 a_n5142_10515.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X327 a_n8898_687.t1 a_n5142_687.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X328 avss.t257 avss.t258 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X329 avss.t228 avss.t229 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X330 a_n15874_4089.t1 a_n12654_3711.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X331 multiplexer_0.trans_gate_m_19.in.t0 multiplexer_0.vtrip_0.t17 multiplexer_0.in_1110.t0 avdd.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X332 avss.t141 multiplexer_0.vtrip_2_b.t6 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X333 comp_hyst_0.net4.t4 comp_hyst_0.net4.t3 dvdd.t8 dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X334 a_n8898_n825.t0 a_n5142_n825.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X335 comp_hyst_0.net3.t8 ena.t7 dvdd.t119 dvdd.t118 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X336 a_n12118_13539.t0 a_n8898_13161.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X337 a_n12654_1065.t1 a_n8898_1065.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X338 avss.t204 avss.t205 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X339 multiplexer_0.trans_gate_m_31.out.t2 multiplexer_0.vtrip_1_b.t10 multiplexer_0.trans_gate_m_31.in.t5 avss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X340 multiplexer_0.trans_gate_m_37.in.t4 multiplexer_0.vtrip_1_b.t11 multiplexer_0.trans_gate_m_18.in.t5 avss.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X341 multiplexer_0.in_0100.t2 multiplexer_0.in_0011.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X342 avss.t153 avss.t154 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X343 comp_hyst_0.net3.t2 comp_hyst_0.net4.t13 dvdd.t7 dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
X344 avss.t102 avss.t103 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X345 a_n15874_7869.t0 a_n12654_7491.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X346 avss.t129 avss.t130 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X347 dvss.t58 dvss.t56 dvss.t57 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X348 a_n15874_n1959.t1 a_n12654_n1581.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X349 a_n8362_10137.t0 a_n5142_10515.t0 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X350 dvss.t3 vtrip[0].t2 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
X351 multiplexer_0.trans_gate_m_33.in.t0 multiplexer_0.vtrip_2_b.t7 multiplexer_0.trans_gate_m_28.in.t0 avdd.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X352 avss.t147 multiplexer_0.vtrip_0_b.t17 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X353 a_n8898_309.t1 a_n5142_n69.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X354 avss.t134 avss.t135 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X355 a_n12118_4467.t0 a_n8898_4845.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X356 avss.t78 avss.t79 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X357 dvss.t75 comp_hyst_0.net5.t0 comp_hyst_0.net5.t1 dvss.t19 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
X358 a_n15874_1065.t1 a_n12654_1443.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X359 a_n12118_11271.t1 a_n8898_10893.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X360 dvss.t55 dvss.t53 dvss.t54 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X361 avss.t145 avss.t146 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X362 a_n8898_14673.t1 a_n5142_14295.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X363 dvss.t1 comp_hyst_0.net2.t3 ovout.t1 dvss.t0 sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
X364 multiplexer_0.in_1000.t1 multiplexer_0.in_1001.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X365 dvss.t5 vtrip[0].t3 level_shifter_0.in_b.t1 dvss.t4 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X366 dvss.t14 comp_hyst_0.ena_b.t4 ovout.t0 dvss.t13 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X367 avss.t132 avss.t133 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X368 multiplexer_0.trans_gate_m_28.in.t4 multiplexer_0.vtrip_1_b.t12 multiplexer_0.trans_gate_m_25.in.t5 avdd.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X369 avss.t76 avss.t77 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X370 a_n15874_n1203.t1 a_n12654_n1203.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X371 multiplexer_0.trans_gate_m_21.in.t4 multiplexer_0.vtrip_0_b.t18 multiplexer_0.in_1010.t3 avss.t239 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X372 a_n12118_2199.t0 a_n8898_1821.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X373 avss.t86 avss.t87 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X374 avss.t174 avss.t175 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X375 dvss.t52 dvss.t50 dvss.t51 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X376 a_n8362_7869.t0 multiplexer_0.in_0010.t3 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X377 a_n15874_12405.t1 a_n12654_12783.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X378 avss.t252 avss.t253 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X379 avss.t64 avss.t65 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X380 avss.t189 multiplexer_0.vtrip_1.t11 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=515385786,232366 d=515385786,232366
X381 dvdd.t35 dvdd.t33 dvdd.t34 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X382 multiplexer_0.trans_gate_m_25.in.t1 multiplexer_0.vtrip_0.t18 multiplexer_0.in_0110.t3 avdd.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X383 avss.t35 avss.t36 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X384 avss.t39 avss.t40 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X385 dvss.t49 dvss.t47 dvss.t48 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X386 multiplexer_0.trans_gate_m_23.in.t1 multiplexer_0.vtrip_0.t19 multiplexer_0.in_1000.t0 avdd.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X387 a_n8362_11649.t1 a_n5142_11271.t1 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X388 a_n12118_8247.t1 a_n8898_8625.t1 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X389 a_n8898_1443.t1 multiplexer_0.in_1111.t2 avss.t13 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X390 dvss.t46 dvss.t44 dvss.t45 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X391 a_n15874_4845.t0 a_n12654_5223.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X392 multiplexer_0.vtrip_1_b.t1 multiplexer_0.vtrip_1.t12 avdd.t19 avdd.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X393 dvss.t43 dvss.t41 dvss.t42 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X394 a_n12118_5979.t1 a_n8898_5601.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X395 a_n15874_2577.t1 a_n12654_2199.t0 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X396 a_n12654_15051.t0 a_n8898_15051.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X397 dvdd.t32 dvdd.t29 dvdd.t31 dvdd.t30 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X398 multiplexer_0.trans_gate_m_31.in.t0 multiplexer_0.vtrip_0.t20 multiplexer_0.in_0001.t0 avss.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X399 vin.t0 multiplexer_0.vtrip_3_b.t5 multiplexer_0.trans_gate_m_37.out.t2 avdd sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X400 dvss.t40 dvss.t38 dvss.t39 dvss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X401 dvss.t37 dvss.t34 dvss.t36 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=1
X402 ibias.t1 comp_hyst_0.ena_b.t5 comp_hyst_0.net5.t2 dvdd.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=5
X403 a_n15874_9381.t1 a_n12654_9003.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X404 a_n15874_12405.t0 a_n12654_12027.t1 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X405 a_n12654_n1959.t1 a_n8898_n1959.t0 avss.t10 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X406 dvss.t33 dvss.t30 dvss.t32 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0 ps=0 w=1.3 l=1
X407 avss.t37 avss.t38 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X408 multiplexer_0.trans_gate_m_19.in.t4 multiplexer_0.vtrip_0_b.t19 multiplexer_0.in_1111.t3 avdd.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X409 multiplexer_0.trans_gate_m_27.in.t3 multiplexer_0.vtrip_0_b.t20 multiplexer_0.in_0100.t3 avss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
X410 avss.t8 avss.t9 avss.t5 sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X411 avss.t62 avss.t63 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X412 avss.t143 avss.t144 avss.t14 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X413 dvdd.t28 dvdd.t26 dvdd.t27 dvdd.t6 sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=8
X414 avss.t159 avss.t160 avss.t0 sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X415 dvss.t10 vtrip[2].t3 sky130_fd_pr__diode_pw2nd_05v5 perim=2.3e+06 area=3.15e+11
**devattr s=153706620,137952 d=153706620,137952
R0 dvss.n449 dvss.n444 254820
R1 dvss.n95 dvss.n94 34996.5
R2 dvss.n94 dvss.n9 31135.3
R3 dvss.n448 dvss.n447 30031.7
R4 dvss.n449 dvss.n448 23444.7
R5 dvss.n533 dvss.n21 17898.5
R6 dvss.n447 dvss.n444 14868.9
R7 dvss.n510 dvss.n54 13807.4
R8 dvss.n510 dvss.n50 13807.4
R9 dvss.n277 dvss.n49 13807.4
R10 dvss.n513 dvss.n49 13807.4
R11 dvss.n566 dvss.n9 13404.2
R12 dvss.n511 dvss.n51 12416.8
R13 dvss.n512 dvss.n511 12416.8
R14 dvss.n464 dvss.n10 11008.6
R15 dvss.n565 dvss.n10 11008.6
R16 dvss.n566 dvss.n565 11008.6
R17 dvss.n528 dvss.n40 6854.44
R18 dvss.n528 dvss.n41 6854.44
R19 dvss.n73 dvss.n41 6854.44
R20 dvss.n73 dvss.n40 6854.44
R21 dvss.n94 dvss.n93 6401.06
R22 dvss.n450 dvss.n443 4698.47
R23 dvss.t2 dvss.n113 4082.08
R24 dvss.n227 dvss.n114 4040.64
R25 dvss.n114 dvss.n105 4040.64
R26 dvss.n250 dvss.n96 4040.64
R27 dvss.n237 dvss.n96 4040.64
R28 dvss.n305 dvss.n69 3957.38
R29 dvss.n302 dvss.n69 3957.38
R30 dvss.n305 dvss.n70 3957.38
R31 dvss.n302 dvss.n70 3957.38
R32 dvss.n460 dvss.n457 3957.38
R33 dvss.n469 dvss.n457 3957.38
R34 dvss.n460 dvss.n459 3957.38
R35 dvss.n484 dvss.n481 3957.38
R36 dvss.n492 dvss.n481 3957.38
R37 dvss.n484 dvss.n483 3957.38
R38 dvss.n552 dvss.n16 3957.38
R39 dvss.n556 dvss.n16 3957.38
R40 dvss.n552 dvss.n18 3957.38
R41 dvss.n299 dvss.n283 3957.38
R42 dvss.n299 dvss.n297 3957.38
R43 dvss.n520 dvss.n516 3957.38
R44 dvss.n521 dvss.n520 3957.38
R45 dvss.n531 dvss.n37 3957.38
R46 dvss.n37 dvss.n35 3957.38
R47 dvss.n36 dvss.n35 3957.38
R48 dvss.n548 dvss.n5 3957.38
R49 dvss.n548 dvss.n546 3957.38
R50 dvss.n571 dvss.n5 3957.38
R51 dvss.n251 dvss.n95 3484.39
R52 dvss.n309 dvss.n308 3186.08
R53 dvss.n127 dvss.n116 3171.26
R54 dvss.n116 dvss.n115 3171.26
R55 dvss.n240 dvss.n112 3171.26
R56 dvss.n240 dvss.n107 3171.26
R57 dvss.n125 dvss.n117 3171.26
R58 dvss.n117 dvss.n106 3171.26
R59 dvss.n124 dvss.n118 3171.26
R60 dvss.n118 dvss.n101 3171.26
R61 dvss.n239 dvss.n238 3171.26
R62 dvss.n239 dvss.n97 3171.26
R63 dvss.n537 dvss.n27 3052.71
R64 dvss.n537 dvss.n536 3052.71
R65 dvss.n536 dvss.n535 3052.71
R66 dvss.n535 dvss.n27 3052.71
R67 dvss.n550 dvss.n21 2973.47
R68 dvss.n446 dvss.n443 2848.04
R69 dvss.n291 dvss.n283 2566.79
R70 dvss.n291 dvss.n290 2566.79
R71 dvss.n290 dvss.n42 2566.79
R72 dvss.n516 dvss.n42 2566.79
R73 dvss.n297 dvss.n284 2566.79
R74 dvss.n289 dvss.n284 2566.79
R75 dvss.n289 dvss.n43 2566.79
R76 dvss.n521 dvss.n43 2566.79
R77 dvss.n21 dvss.n9 2126.29
R78 dvss.n459 dvss.n455 1836.74
R79 dvss.n483 dvss.n479 1836.74
R80 dvss.n18 dvss.n15 1836.74
R81 dvss.n546 dvss.n3 1836.74
R82 dvss.n84 dvss.n58 1735.47
R83 dvss.n312 dvss.n58 1735.47
R84 dvss.n253 dvss.n92 1735.47
R85 dvss.n187 dvss.n181 1735.47
R86 dvss.n187 dvss.n157 1735.47
R87 dvss.n171 dvss.n170 1735.47
R88 dvss.n465 dvss.n458 1720.85
R89 dvss.n488 dvss.n482 1720.85
R90 dvss.n564 dvss.n11 1720.85
R91 dvss.n567 dvss.n6 1720.85
R92 dvss.t11 dvss.n19 1584.72
R93 dvss.n465 dvss.n456 1552.82
R94 dvss.n472 dvss.n456 1552.82
R95 dvss.n488 dvss.n480 1552.82
R96 dvss.n495 dvss.n480 1552.82
R97 dvss.n564 dvss.n12 1552.82
R98 dvss.n559 dvss.n12 1552.82
R99 dvss.n540 dvss.n22 1552.82
R100 dvss.n544 dvss.n22 1552.82
R101 dvss.n540 dvss.n23 1552.82
R102 dvss.n544 dvss.n23 1552.82
R103 dvss.n149 dvss.n132 1552.82
R104 dvss.n133 dvss.n132 1552.82
R105 dvss.n149 dvss.n148 1552.82
R106 dvss.n148 dvss.n133 1552.82
R107 dvss.n220 dvss.n219 1552.82
R108 dvss.n221 dvss.n220 1552.82
R109 dvss.n222 dvss.n219 1552.82
R110 dvss.n222 dvss.n221 1552.82
R111 dvss.n574 dvss.n4 1552.82
R112 dvss.n567 dvss.n4 1552.82
R113 dvss.n469 dvss.n458 1390.59
R114 dvss.n492 dvss.n482 1390.59
R115 dvss.n556 dvss.n11 1390.59
R116 dvss.n525 dvss.n42 1390.59
R117 dvss.n525 dvss.n43 1390.59
R118 dvss.n292 dvss.n291 1390.59
R119 dvss.n292 dvss.n284 1390.59
R120 dvss.n54 dvss.n51 1390.59
R121 dvss.n277 dvss.n51 1390.59
R122 dvss.n513 dvss.n512 1390.59
R123 dvss.n512 dvss.n50 1390.59
R124 dvss.n571 dvss.n6 1390.59
R125 dvss.t21 dvss.n20 1254.31
R126 dvss.n551 dvss.t8 1254.31
R127 dvss.n549 dvss.t4 1254.31
R128 dvss.n471 dvss.t11 1133.98
R129 dvss.n169 dvss.t31 1114.84
R130 dvss.n252 dvss.t35 1114.84
R131 dvss.n271 dvss.n60 968.173
R132 dvss.n60 dvss.n57 968.173
R133 dvss.n259 dvss.n79 968.173
R134 dvss.n270 dvss.n79 968.173
R135 dvss.n270 dvss.n269 968.173
R136 dvss.n269 dvss.n80 968.173
R137 dvss.n64 dvss.n59 968.173
R138 dvss.n260 dvss.n59 968.173
R139 dvss.n260 dvss.n62 968.173
R140 dvss.n271 dvss.n62 968.173
R141 dvss.n267 dvss.n85 968.173
R142 dvss.n267 dvss.n87 968.173
R143 dvss.n87 dvss.n82 968.173
R144 dvss.n259 dvss.n82 968.173
R145 dvss.n310 dvss.n63 968.173
R146 dvss.n310 dvss.n64 968.173
R147 dvss.n107 dvss.n104 968.173
R148 dvss.n115 dvss.n104 968.173
R149 dvss.n229 dvss.n125 968.173
R150 dvss.n229 dvss.n112 968.173
R151 dvss.n126 dvss.n112 968.173
R152 dvss.n127 dvss.n126 968.173
R153 dvss.n103 dvss.n101 968.173
R154 dvss.n106 dvss.n103 968.173
R155 dvss.n244 dvss.n106 968.173
R156 dvss.n244 dvss.n107 968.173
R157 dvss.n238 dvss.n120 968.173
R158 dvss.n124 dvss.n120 968.173
R159 dvss.n231 dvss.n124 968.173
R160 dvss.n231 dvss.n125 968.173
R161 dvss.n246 dvss.n97 968.173
R162 dvss.n246 dvss.n101 968.173
R163 dvss.n203 dvss.n156 968.173
R164 dvss.n192 dvss.n156 968.173
R165 dvss.n208 dvss.n178 968.173
R166 dvss.n208 dvss.n182 968.173
R167 dvss.n182 dvss.n180 968.173
R168 dvss.n191 dvss.n180 968.173
R169 dvss.n160 dvss.n155 968.173
R170 dvss.n197 dvss.n155 968.173
R171 dvss.n197 dvss.n158 968.173
R172 dvss.n203 dvss.n158 968.173
R173 dvss.n177 dvss.n164 968.173
R174 dvss.n211 dvss.n177 968.173
R175 dvss.n211 dvss.n210 968.173
R176 dvss.n210 dvss.n178 968.173
R177 dvss.n216 dvss.n159 968.173
R178 dvss.n216 dvss.n160 968.173
R179 dvss.n494 dvss.t21 897.556
R180 dvss.n558 dvss.t8 897.556
R181 dvss.n573 dvss.t4 897.556
R182 dvss.n84 dvss.n80 869.38
R183 dvss.n312 dvss.n57 869.38
R184 dvss.n90 dvss.n63 869.38
R185 dvss.n253 dvss.n85 869.38
R186 dvss.n227 dvss.n127 869.38
R187 dvss.n115 dvss.n105 869.38
R188 dvss.n250 dvss.n97 869.38
R189 dvss.n238 dvss.n237 869.38
R190 dvss.n191 dvss.n181 869.38
R191 dvss.n192 dvss.n157 869.38
R192 dvss.n170 dvss.n159 869.38
R193 dvss.n173 dvss.n164 869.38
R194 dvss.n139 dvss.n80 866.087
R195 dvss.n139 dvss.n57 866.087
R196 dvss.n272 dvss.n270 866.087
R197 dvss.n272 dvss.n271 866.087
R198 dvss.n261 dvss.n259 866.087
R199 dvss.n261 dvss.n260 866.087
R200 dvss.n87 dvss.n86 866.087
R201 dvss.n86 dvss.n64 866.087
R202 dvss.n255 dvss.n85 866.087
R203 dvss.n255 dvss.n63 866.087
R204 dvss.n193 dvss.n191 866.087
R205 dvss.n193 dvss.n192 866.087
R206 dvss.n204 dvss.n182 866.087
R207 dvss.n204 dvss.n203 866.087
R208 dvss.n198 dvss.n178 866.087
R209 dvss.n198 dvss.n197 866.087
R210 dvss.n212 dvss.n211 866.087
R211 dvss.n212 dvss.n160 866.087
R212 dvss.n165 dvss.n164 866.087
R213 dvss.n165 dvss.n159 866.087
R214 dvss.n275 dvss.n52 800.378
R215 dvss.n52 dvss.n48 800.378
R216 dvss.n458 dvss.n455 730.059
R217 dvss.n482 dvss.n479 730.059
R218 dvss.n15 dvss.n11 730.059
R219 dvss.n6 dvss.n3 730.059
R220 dvss.n91 dvss.n90 686.495
R221 dvss.n173 dvss.n172 686.495
R222 dvss.n472 dvss.n455 654.736
R223 dvss.n495 dvss.n479 654.736
R224 dvss.n559 dvss.n15 654.736
R225 dvss.n574 dvss.n3 654.736
R226 dvss.n543 dvss.n542 627.953
R227 dvss.n464 dvss.t17 543.74
R228 dvss.n169 dvss.n113 474.76
R229 dvss.n252 dvss.n251 474.76
R230 dvss.n249 dvss.n98 466.447
R231 dvss.n236 dvss.n98 466.447
R232 dvss.n471 dvss.n470 450.733
R233 dvss.n74 dvss.n72 445.365
R234 dvss.t10 dvss.n10 430.373
R235 dvss.n565 dvss.t7 430.373
R236 dvss.n566 dvss.t3 430.373
R237 dvss.n542 dvss.n541 429.183
R238 dvss.t2 dvss.n119 396.166
R239 dvss.n534 dvss.t29 374.048
R240 dvss.n538 dvss.t29 374.048
R241 dvss.n235 dvss.n99 362.541
R242 dvss.n248 dvss.n99 362.541
R243 dvss.n233 dvss.n121 362.541
R244 dvss.n121 dvss.n100 362.541
R245 dvss.n123 dvss.n122 362.541
R246 dvss.n122 dvss.n109 362.541
R247 dvss.n241 dvss.n111 362.541
R248 dvss.n242 dvss.n241 362.541
R249 dvss.n134 dvss.n129 362.541
R250 dvss.n135 dvss.n134 362.541
R251 dvss.n494 dvss.n493 356.757
R252 dvss.n558 dvss.n557 356.757
R253 dvss.n573 dvss.n572 356.757
R254 dvss.n30 dvss.n29 353.507
R255 dvss.n72 dvss.n38 348.613
R256 dvss.n102 dvss.n95 331.055
R257 dvss.n451 dvss.n442 305.281
R258 dvss.n465 dvss.n464 303.233
R259 dvss.n488 dvss.n10 300.995
R260 dvss.n565 dvss.n564 300.995
R261 dvss.n567 dvss.n566 300.995
R262 dvss.n542 dvss.n23 293.281
R263 dvss.n466 dvss.n465 292.5
R264 dvss.n463 dvss.n456 292.5
R265 dvss.t17 dvss.n456 292.5
R266 dvss.n473 dvss.n472 292.5
R267 dvss.n472 dvss.n471 292.5
R268 dvss.n489 dvss.n488 292.5
R269 dvss.n487 dvss.n480 292.5
R270 dvss.t10 dvss.n480 292.5
R271 dvss.n496 dvss.n495 292.5
R272 dvss.n495 dvss.n494 292.5
R273 dvss.n564 dvss.n563 292.5
R274 dvss.n562 dvss.n12 292.5
R275 dvss.n12 dvss.t7 292.5
R276 dvss.n560 dvss.n559 292.5
R277 dvss.n559 dvss.n558 292.5
R278 dvss.n221 dvss.n152 292.5
R279 dvss.n221 dvss.n119 292.5
R280 dvss.n223 dvss.n222 292.5
R281 dvss.n222 dvss.t6 292.5
R282 dvss.n219 dvss.n154 292.5
R283 dvss.n219 dvss.n218 292.5
R284 dvss.n220 dvss.n130 292.5
R285 dvss.n220 dvss.t6 292.5
R286 dvss.n145 dvss.n133 292.5
R287 dvss.n133 dvss.n83 292.5
R288 dvss.n148 dvss.n147 292.5
R289 dvss.n148 dvss.t18 292.5
R290 dvss.n150 dvss.n149 292.5
R291 dvss.n149 dvss.n102 292.5
R292 dvss.n138 dvss.n132 292.5
R293 dvss.n132 dvss.t18 292.5
R294 dvss.n544 dvss.n543 292.5
R295 dvss.n545 dvss.n544 292.5
R296 dvss.n23 dvss.t74 292.5
R297 dvss.n541 dvss.n540 292.5
R298 dvss.n540 dvss.n539 292.5
R299 dvss.n24 dvss.n22 292.5
R300 dvss.n22 dvss.t74 292.5
R301 dvss.n8 dvss.n4 292.5
R302 dvss.t3 dvss.n4 292.5
R303 dvss.n568 dvss.n567 292.5
R304 dvss.n575 dvss.n574 292.5
R305 dvss.n574 dvss.n573 292.5
R306 dvss.n515 dvss.n47 292.142
R307 dvss.n515 dvss.n514 292.142
R308 dvss.n462 dvss.n461 257.13
R309 dvss.n486 dvss.n485 257.13
R310 dvss.n554 dvss.n553 257.13
R311 dvss.n47 dvss.n46 257.13
R312 dvss.n547 dvss.n7 257.13
R313 dvss.n29 dvss.n28 246.004
R314 dvss.n570 dvss.n7 215.569
R315 dvss.n303 dvss.n71 215.506
R316 dvss.n533 dvss.t27 215.23
R317 dvss.n298 dvss.t13 203.126
R318 dvss.t25 dvss.n53 203.126
R319 dvss.n526 dvss.t23 203.126
R320 dvss.n89 dvss.n88 202.918
R321 dvss.n254 dvss.n88 202.918
R322 dvss.n168 dvss.n167 202.918
R323 dvss.n174 dvss.n167 202.918
R324 dvss.n533 dvss.n31 192.123
R325 dvss.n550 dvss.n19 189.595
R326 dvss.n445 dvss.n442 185.155
R327 dvss.n468 dvss.n462 175.536
R328 dvss.n491 dvss.n486 175.536
R329 dvss.n555 dvss.n554 175.536
R330 dvss.t13 dvss.t15 173.322
R331 dvss.n46 dvss.n38 169.59
R332 dvss.t27 dvss.t23 160.484
R333 dvss.n33 dvss.n31 160.484
R334 dvss.n311 dvss.n61 150.856
R335 dvss.n550 dvss.n20 150.065
R336 dvss.n551 dvss.n550 150.065
R337 dvss.n550 dvss.n549 150.065
R338 dvss.n316 dvss.n30 148.329
R339 dvss.n527 dvss.n34 146.728
R340 dvss.n550 dvss.n545 129.994
R341 dvss.n315 dvss.n50 126.078
R342 dvss.n414 dvss.t44 125.236
R343 dvss.t44 dvss.n413 125.236
R344 dvss.n394 dvss.t68 125.236
R345 dvss.t68 dvss.n393 125.236
R346 dvss.n390 dvss.t71 125.236
R347 dvss.t71 dvss.n389 125.236
R348 dvss.n386 dvss.t41 125.236
R349 dvss.t41 dvss.n385 125.236
R350 dvss.n382 dvss.t30 125.236
R351 dvss.t30 dvss.n381 125.236
R352 dvss.t47 dvss.n417 125.236
R353 dvss.n418 dvss.t47 125.236
R354 dvss.n323 dvss.t53 125.236
R355 dvss.t53 dvss.n322 125.236
R356 dvss.n321 dvss.t50 125.236
R357 dvss.t50 dvss.n320 125.236
R358 dvss.n445 dvss.n444 122.587
R359 dvss.n209 dvss.t31 120.593
R360 dvss.n311 dvss.t35 120.593
R361 dvss.n316 dvss.n25 120.013
R362 dvss.n373 dvss.t59 118.005
R363 dvss.t59 dvss.n372 118.005
R364 dvss.n360 dvss.t56 118.005
R365 dvss.t56 dvss.n355 118.005
R366 dvss.n410 dvss.t34 118.005
R367 dvss.t34 dvss.n409 118.005
R368 dvss.n400 dvss.t65 118.005
R369 dvss.t65 dvss.n399 118.005
R370 dvss.n469 dvss.n468 117.001
R371 dvss.n470 dvss.n469 117.001
R372 dvss.n461 dvss.n460 117.001
R373 dvss.n460 dvss.n19 117.001
R374 dvss.n492 dvss.n491 117.001
R375 dvss.n493 dvss.n492 117.001
R376 dvss.n485 dvss.n484 117.001
R377 dvss.n484 dvss.n20 117.001
R378 dvss.n556 dvss.n555 117.001
R379 dvss.n557 dvss.n556 117.001
R380 dvss.n553 dvss.n552 117.001
R381 dvss.n552 dvss.n551 117.001
R382 dvss.n171 dvss.n167 117.001
R383 dvss.n166 dvss.n165 117.001
R384 dvss.n165 dvss.t31 117.001
R385 dvss.n92 dvss.n88 117.001
R386 dvss.n256 dvss.n255 117.001
R387 dvss.n255 dvss.t35 117.001
R388 dvss.n47 dvss.n35 117.001
R389 dvss.t27 dvss.n35 117.001
R390 dvss.n531 dvss.n530 117.001
R391 dvss.n213 dvss.n212 117.001
R392 dvss.n212 dvss.t31 117.001
R393 dvss.n199 dvss.n198 117.001
R394 dvss.n198 dvss.t31 117.001
R395 dvss.n205 dvss.n204 117.001
R396 dvss.n204 dvss.t31 117.001
R397 dvss.n194 dvss.n193 117.001
R398 dvss.n193 dvss.t31 117.001
R399 dvss.n188 dvss.n187 117.001
R400 dvss.n187 dvss.t31 117.001
R401 dvss.n514 dvss.n513 117.001
R402 dvss.n513 dvss.n31 117.001
R403 dvss.n50 dvss.n31 117.001
R404 dvss.n55 dvss.n54 117.001
R405 dvss.n61 dvss.n54 117.001
R406 dvss.n278 dvss.n277 117.001
R407 dvss.n277 dvss.n61 117.001
R408 dvss.n293 dvss.n292 117.001
R409 dvss.n292 dvss.n53 117.001
R410 dvss.n525 dvss.n524 117.001
R411 dvss.n526 dvss.n525 117.001
R412 dvss.n520 dvss.n519 117.001
R413 dvss.n520 dvss.n33 117.001
R414 dvss.n300 dvss.n299 117.001
R415 dvss.n299 dvss.n298 117.001
R416 dvss.n281 dvss.n70 117.001
R417 dvss.t0 dvss.n70 117.001
R418 dvss.n69 dvss.n66 117.001
R419 dvss.t0 dvss.n69 117.001
R420 dvss.n529 dvss.n528 117.001
R421 dvss.n528 dvss.n527 117.001
R422 dvss.n74 dvss.n73 117.001
R423 dvss.n73 dvss.n71 117.001
R424 dvss.n86 dvss.n67 117.001
R425 dvss.n86 dvss.t35 117.001
R426 dvss.n262 dvss.n261 117.001
R427 dvss.n261 dvss.t35 117.001
R428 dvss.n273 dvss.n272 117.001
R429 dvss.n272 dvss.t35 117.001
R430 dvss.n140 dvss.n139 117.001
R431 dvss.n139 dvss.t35 117.001
R432 dvss.n144 dvss.n58 117.001
R433 dvss.t35 dvss.n58 117.001
R434 dvss.n571 dvss.n570 117.001
R435 dvss.n572 dvss.n571 117.001
R436 dvss.n548 dvss.n547 117.001
R437 dvss.n549 dvss.n548 117.001
R438 dvss.n235 dvss.n234 115.201
R439 dvss.n234 dvss.n233 115.201
R440 dvss.n248 dvss.n247 115.201
R441 dvss.n247 dvss.n100 115.201
R442 dvss.n108 dvss.n100 115.201
R443 dvss.n109 dvss.n108 115.201
R444 dvss.n233 dvss.n232 115.201
R445 dvss.n232 dvss.n123 115.201
R446 dvss.n228 dvss.n123 115.201
R447 dvss.n228 dvss.n111 115.201
R448 dvss.n243 dvss.n109 115.201
R449 dvss.n243 dvss.n242 115.201
R450 dvss.n242 dvss.n110 115.201
R451 dvss.n135 dvss.n110 115.201
R452 dvss.n128 dvss.n111 115.201
R453 dvss.n129 dvss.n128 115.201
R454 dvss.n81 dvss.n78 115.201
R455 dvss.n141 dvss.n81 115.201
R456 dvss.n263 dvss.n258 115.201
R457 dvss.n258 dvss.n78 115.201
R458 dvss.n265 dvss.n264 115.201
R459 dvss.n264 dvss.n263 115.201
R460 dvss.n266 dvss.n257 115.201
R461 dvss.n266 dvss.n265 115.201
R462 dvss.n309 dvss.n65 115.201
R463 dvss.n202 dvss.n196 115.201
R464 dvss.n196 dvss.n195 115.201
R465 dvss.n207 dvss.n183 115.201
R466 dvss.n207 dvss.n206 115.201
R467 dvss.n206 dvss.n184 115.201
R468 dvss.n190 dvss.n184 115.201
R469 dvss.n214 dvss.n162 115.201
R470 dvss.n200 dvss.n162 115.201
R471 dvss.n201 dvss.n200 115.201
R472 dvss.n202 dvss.n201 115.201
R473 dvss.n176 dvss.n175 115.201
R474 dvss.n176 dvss.n163 115.201
R475 dvss.n179 dvss.n163 115.201
R476 dvss.n183 dvss.n179 115.201
R477 dvss.n215 dvss.n161 115.201
R478 dvss.n215 dvss.n214 115.201
R479 dvss.n189 dvss.n188 112.451
R480 dvss.n532 dvss.n531 112.177
R481 dvss.n304 dvss.t0 111.421
R482 dvss.t0 dvss.n303 111.421
R483 dvss.n75 dvss.n66 104.514
R484 dvss.n249 dvss.n248 103.906
R485 dvss.n236 dvss.n235 103.906
R486 dvss.n226 dvss.n129 103.906
R487 dvss.n226 dvss.n225 103.906
R488 dvss.n136 dvss.n135 103.906
R489 dvss.n137 dvss.n136 103.906
R490 dvss.n142 dvss.n141 103.906
R491 dvss.n143 dvss.n142 103.906
R492 dvss.n89 dvss.n65 103.906
R493 dvss.n257 dvss.n254 103.906
R494 dvss.n190 dvss.n189 103.906
R495 dvss.n195 dvss.n186 103.906
R496 dvss.n186 dvss.n185 103.906
R497 dvss.n168 dvss.n161 103.906
R498 dvss.n175 dvss.n174 103.906
R499 dvss.n470 dvss.t17 103.74
R500 dvss.n461 dvss.n453 100.233
R501 dvss.n485 dvss.n477 100.233
R502 dvss.n553 dvss.n17 100.233
R503 dvss.n547 dvss.n1 100.233
R504 dvss.n141 dvss.n140 99.0123
R505 dvss.n273 dvss.n78 99.0123
R506 dvss.n263 dvss.n262 99.0123
R507 dvss.n265 dvss.n67 99.0123
R508 dvss.n257 dvss.n256 99.0123
R509 dvss.n256 dvss.n65 99.0123
R510 dvss.n194 dvss.n190 99.0123
R511 dvss.n195 dvss.n194 99.0123
R512 dvss.n206 dvss.n205 99.0123
R513 dvss.n205 dvss.n202 99.0123
R514 dvss.n199 dvss.n183 99.0123
R515 dvss.n200 dvss.n199 99.0123
R516 dvss.n213 dvss.n163 99.0123
R517 dvss.n214 dvss.n213 99.0123
R518 dvss.n175 dvss.n166 99.0123
R519 dvss.n166 dvss.n161 99.0123
R520 dvss.n174 dvss.n173 97.5005
R521 dvss.n170 dvss.n168 97.5005
R522 dvss.n170 dvss.n169 97.5005
R523 dvss.n237 dvss.n236 97.5005
R524 dvss.n237 dvss.n113 97.5005
R525 dvss.n250 dvss.n249 97.5005
R526 dvss.n251 dvss.n250 97.5005
R527 dvss.n254 dvss.n253 97.5005
R528 dvss.n253 dvss.n252 97.5005
R529 dvss.n90 dvss.n89 97.5005
R530 dvss.n189 dvss.n181 97.5005
R531 dvss.n209 dvss.n181 97.5005
R532 dvss.n186 dvss.n157 97.5005
R533 dvss.n217 dvss.n157 97.5005
R534 dvss.n227 dvss.n226 97.5005
R535 dvss.n230 dvss.n227 97.5005
R536 dvss.n136 dvss.n105 97.5005
R537 dvss.n245 dvss.n105 97.5005
R538 dvss.n142 dvss.n84 97.5005
R539 dvss.n268 dvss.n84 97.5005
R540 dvss.n313 dvss.n312 97.5005
R541 dvss.n312 dvss.n311 97.5005
R542 dvss.n535 dvss.n30 97.5005
R543 dvss.n535 dvss.n534 97.5005
R544 dvss.n537 dvss.n26 97.5005
R545 dvss.n538 dvss.n537 97.5005
R546 dvss.n514 dvss.n48 96.7534
R547 dvss.n524 dvss.n44 94.3698
R548 dvss.n140 dvss.n56 92.6123
R549 dvss.n276 dvss.n273 92.6123
R550 dvss.n262 dvss.n77 92.6123
R551 dvss.n307 dvss.n67 92.6123
R552 dvss.n304 dvss.n61 91.7054
R553 dvss.n524 dvss.n523 90.3534
R554 dvss.n293 dvss.n287 90.3534
R555 dvss.n294 dvss.n293 90.3534
R556 dvss.n308 dvss.n66 85.0829
R557 dvss.n423 dvss.t28 84.6474
R558 dvss.n422 dvss.t16 84.2828
R559 dvss.n476 dvss.t12 84.2462
R560 dvss.n499 dvss.t22 84.2462
R561 dvss.n501 dvss.t9 84.2462
R562 dvss.n0 dvss.t5 84.2462
R563 dvss.n318 dvss.t20 83.7172
R564 dvss.n429 dvss.t75 83.7172
R565 dvss.n420 dvss.t14 83.7172
R566 dvss.n425 dvss.t26 83.7172
R567 dvss.n421 dvss.t24 83.7172
R568 dvss.n177 dvss.n176 83.5719
R569 dvss.n209 dvss.n177 83.5719
R570 dvss.n216 dvss.n215 83.5719
R571 dvss.n217 dvss.n216 83.5719
R572 dvss.n210 dvss.n179 83.5719
R573 dvss.n210 dvss.n209 83.5719
R574 dvss.n162 dvss.n155 83.5719
R575 dvss.n217 dvss.n155 83.5719
R576 dvss.n208 dvss.n207 83.5719
R577 dvss.n209 dvss.n208 83.5719
R578 dvss.n201 dvss.n158 83.5719
R579 dvss.n217 dvss.n158 83.5719
R580 dvss.n184 dvss.n180 83.5719
R581 dvss.n209 dvss.n180 83.5719
R582 dvss.n196 dvss.n156 83.5719
R583 dvss.n217 dvss.n156 83.5719
R584 dvss.n234 dvss.n120 83.5719
R585 dvss.n230 dvss.n120 83.5719
R586 dvss.n247 dvss.n246 83.5719
R587 dvss.n246 dvss.n245 83.5719
R588 dvss.n232 dvss.n231 83.5719
R589 dvss.n231 dvss.n230 83.5719
R590 dvss.n108 dvss.n103 83.5719
R591 dvss.n245 dvss.n103 83.5719
R592 dvss.n229 dvss.n228 83.5719
R593 dvss.n230 dvss.n229 83.5719
R594 dvss.n244 dvss.n243 83.5719
R595 dvss.n245 dvss.n244 83.5719
R596 dvss.n128 dvss.n126 83.5719
R597 dvss.n230 dvss.n126 83.5719
R598 dvss.n110 dvss.n104 83.5719
R599 dvss.n245 dvss.n104 83.5719
R600 dvss.n267 dvss.n266 83.5719
R601 dvss.n268 dvss.n267 83.5719
R602 dvss.n310 dvss.n309 83.5719
R603 dvss.n311 dvss.n310 83.5719
R604 dvss.n264 dvss.n82 83.5719
R605 dvss.n268 dvss.n82 83.5719
R606 dvss.n68 dvss.n59 83.5719
R607 dvss.n311 dvss.n59 83.5719
R608 dvss.n258 dvss.n79 83.5719
R609 dvss.n268 dvss.n79 83.5719
R610 dvss.n279 dvss.n62 83.5719
R611 dvss.n311 dvss.n62 83.5719
R612 dvss.n269 dvss.n81 83.5719
R613 dvss.n269 dvss.n268 83.5719
R614 dvss.n274 dvss.n60 83.5719
R615 dvss.n311 dvss.n60 83.5719
R616 dvss.n438 dvss.t61 82.8472
R617 dvss.n359 dvss.t57 82.8472
R618 dvss.n354 dvss.t58 82.8472
R619 dvss.n364 dvss.t60 82.8472
R620 dvss.n407 dvss.t36 82.8472
R621 dvss.n397 dvss.t66 82.8472
R622 dvss.n332 dvss.t37 82.8472
R623 dvss.n334 dvss.t64 82.8472
R624 dvss.n336 dvss.t63 82.8472
R625 dvss.n338 dvss.t67 82.8472
R626 dvss.n363 dvss.t40 82.8472
R627 dvss.n356 dvss.t39 82.8472
R628 dvss.n493 dvss.t10 82.1112
R629 dvss.n557 dvss.t7 82.1112
R630 dvss.n572 dvss.t3 82.1112
R631 dvss.n433 dvss.t55 77.4826
R632 dvss.n436 dvss.t52 77.4826
R633 dvss.n369 dvss.t51 77.4826
R634 dvss.n366 dvss.t54 77.4826
R635 dvss.n326 dvss.t48 77.4826
R636 dvss.n324 dvss.t49 77.4826
R637 dvss.n330 dvss.t45 77.4826
R638 dvss.n328 dvss.t46 77.4826
R639 dvss.n339 dvss.t69 77.4826
R640 dvss.n344 dvss.t72 77.4826
R641 dvss.n348 dvss.t42 77.4826
R642 dvss.n352 dvss.t32 77.4826
R643 dvss.n350 dvss.t33 77.4826
R644 dvss.n346 dvss.t43 77.4826
R645 dvss.n342 dvss.t73 77.4826
R646 dvss.n341 dvss.t70 77.4826
R647 dvss.n569 dvss.n568 77.3462
R648 dvss.n569 dvss.n2 75.6711
R649 dvss.n83 dvss.t35 75.657
R650 dvss.n218 dvss.t31 75.1985
R651 dvss.n539 dvss.t74 73.3432
R652 dvss.n545 dvss.t74 73.3432
R653 dvss.n172 dvss.n171 66.2531
R654 dvss.n92 dvss.n91 66.2531
R655 dvss.t2 dvss.n95 58.3417
R656 dvss.n543 dvss.n24 57.3914
R657 dvss.n539 dvss.n538 56.418
R658 dvss.n298 dvss.n71 55.9405
R659 dvss.n534 dvss.n533 55.2896
R660 dvss.n459 dvss.n453 53.1823
R661 dvss.n459 dvss.t11 53.1823
R662 dvss.n462 dvss.n457 53.1823
R663 dvss.n457 dvss.t11 53.1823
R664 dvss.n483 dvss.n477 53.1823
R665 dvss.n483 dvss.t21 53.1823
R666 dvss.n486 dvss.n481 53.1823
R667 dvss.n481 dvss.t21 53.1823
R668 dvss.n18 dvss.n17 53.1823
R669 dvss.n18 dvss.t8 53.1823
R670 dvss.n554 dvss.n16 53.1823
R671 dvss.n16 dvss.t8 53.1823
R672 dvss.n46 dvss.n37 53.1823
R673 dvss.n93 dvss.n37 53.1823
R674 dvss.n522 dvss.n521 53.1823
R675 dvss.n521 dvss.t23 53.1823
R676 dvss.n289 dvss.n45 53.1823
R677 dvss.t25 dvss.n289 53.1823
R678 dvss.n297 dvss.n296 53.1823
R679 dvss.t13 dvss.n297 53.1823
R680 dvss.n285 dvss.n283 53.1823
R681 dvss.t13 dvss.n283 53.1823
R682 dvss.n290 dvss.n288 53.1823
R683 dvss.n290 dvss.t25 53.1823
R684 dvss.n517 dvss.n516 53.1823
R685 dvss.n516 dvss.t23 53.1823
R686 dvss.n302 dvss.n301 53.1823
R687 dvss.n303 dvss.n302 53.1823
R688 dvss.n306 dvss.n305 53.1823
R689 dvss.n305 dvss.n304 53.1823
R690 dvss.n518 dvss.n36 53.1823
R691 dvss.n7 dvss.n5 53.1823
R692 dvss.n5 dvss.t4 53.1823
R693 dvss.n546 dvss.n1 53.1823
R694 dvss.n546 dvss.t4 53.1823
R695 dvss.t25 dvss.n34 52.7308
R696 dvss.n147 dvss.n131 51.9534
R697 dvss.n147 dvss.n146 51.9534
R698 dvss.n223 dvss.n153 51.9534
R699 dvss.n224 dvss.n223 51.9534
R700 dvss.n532 dvss.n36 50.9901
R701 dvss.n466 dvss.n463 49.0248
R702 dvss.n489 dvss.n487 49.0248
R703 dvss.n563 dvss.n562 49.0248
R704 dvss.n568 dvss.n8 49.0248
R705 dvss.n172 dvss.t31 46.2824
R706 dvss.n91 dvss.t35 46.2824
R707 dvss.n75 dvss.n74 45.9798
R708 dvss.n245 dvss.n102 45.8529
R709 dvss.n218 dvss.n217 45.3944
R710 dvss.n230 dvss.n119 45.3944
R711 dvss.n268 dvss.n83 44.9359
R712 dvss.n93 dvss.n32 44.3777
R713 dvss.n467 dvss.n466 43.6573
R714 dvss.n490 dvss.n489 43.6573
R715 dvss.n563 dvss.n13 43.6573
R716 dvss.t27 dvss.n33 42.6433
R717 dvss.t15 dvss.n34 37.7211
R718 dvss.n315 dvss.n48 36.3262
R719 dvss.n467 dvss.n454 34.6358
R720 dvss.n490 dvss.n478 34.6358
R721 dvss.n561 dvss.n13 34.6358
R722 dvss.n29 dvss.n27 34.4123
R723 dvss.n27 dvss.t29 34.4123
R724 dvss.n536 dvss.n25 34.4123
R725 dvss.n536 dvss.t29 34.4123
R726 dvss.n522 dvss.n515 31.827
R727 dvss.n428 dvss.t1 30.767
R728 dvss.n509 dvss.n314 29.5006
R729 dvss.n152 dvss.n151 28.0695
R730 dvss.n151 dvss.n150 28.037
R731 dvss.n268 dvss.t18 26.1364
R732 dvss.n217 dvss.t6 25.6779
R733 dvss.n230 dvss.t6 25.6779
R734 dvss.n533 dvss.n32 25.5174
R735 dvss.n245 dvss.t18 25.2193
R736 dvss.n72 dvss.n40 23.4005
R737 dvss.n40 dvss.n32 23.4005
R738 dvss.n286 dvss.n41 23.4005
R739 dvss.t15 dvss.n41 23.4005
R740 dvss.n288 dvss.n287 23.0509
R741 dvss.n98 dvss.n96 22.5005
R742 dvss.t2 dvss.n96 22.5005
R743 dvss.n239 dvss.n99 22.5005
R744 dvss.t2 dvss.n239 22.5005
R745 dvss.n121 dvss.n118 22.5005
R746 dvss.t2 dvss.n118 22.5005
R747 dvss.n122 dvss.n117 22.5005
R748 dvss.t2 dvss.n117 22.5005
R749 dvss.n241 dvss.n240 22.5005
R750 dvss.n240 dvss.t2 22.5005
R751 dvss.n134 dvss.n116 22.5005
R752 dvss.t2 dvss.n116 22.5005
R753 dvss.n151 dvss.n114 22.5005
R754 dvss.t2 dvss.n114 22.5005
R755 dvss.n285 dvss.n76 22.1664
R756 dvss.n288 dvss.n44 21.7501
R757 dvss.n452 dvss.n451 21.6109
R758 dvss.t19 dvss.t15 20.1756
R759 dvss.n286 dvss.n285 19.6688
R760 dvss.n294 dvss.n45 18.5312
R761 dvss.n523 dvss.n45 18.5312
R762 dvss.n523 dvss.n522 18.5312
R763 dvss.n508 dvss.n317 18.0964
R764 dvss.n296 dvss.n282 17.8201
R765 dvss.n296 dvss.n295 17.6528
R766 dvss.n519 dvss.n518 17.4088
R767 dvss.n518 dvss.n517 15.6648
R768 dvss.n468 dvss.n467 15.1599
R769 dvss.n491 dvss.n490 15.1599
R770 dvss.n555 dvss.n13 15.1599
R771 dvss.n317 dvss.n315 14.2671
R772 dvss.n570 dvss.n569 14.1572
R773 dvss.n509 dvss.n508 13.7723
R774 dvss.n542 dvss.n25 13.1595
R775 dvss.n541 dvss.n26 12.8005
R776 dvss.t38 dvss.n376 11.7013
R777 dvss.n377 dvss.t38 11.7013
R778 dvss.t62 dvss.n404 11.7013
R779 dvss.n405 dvss.t62 11.7013
R780 dvss.n529 dvss.n39 11.2005
R781 dvss.n282 dvss.n281 10.4113
R782 dvss.n281 dvss.n280 10.1864
R783 dvss.t19 dvss.n53 9.62951
R784 dvss.n511 dvss.n52 9.59066
R785 dvss.n511 dvss.t19 9.59066
R786 dvss.n510 dvss.n509 9.59066
R787 dvss.t19 dvss.n510 9.59066
R788 dvss.n295 dvss.n49 9.59066
R789 dvss.t19 dvss.n49 9.59066
R790 dvss.n314 dvss.n55 8.46331
R791 dvss.n300 dvss.n282 8.03628
R792 dvss.n144 dvss.n56 7.99238
R793 dvss.n137 dvss.n131 7.92886
R794 dvss.n225 dvss.n224 7.83334
R795 dvss.n185 dvss.n153 7.83334
R796 dvss.n146 dvss.n143 7.73781
R797 dvss.n28 dvss.n24 7.52991
R798 dvss.n275 dvss.n274 7.47598
R799 dvss.n77 dvss.n68 7.34402
R800 dvss.n530 dvss.n38 7.08621
R801 dvss.n143 dvss.n138 6.74438
R802 dvss.t27 dvss.n34 6.65708
R803 dvss.n185 dvss.n130 6.61638
R804 dvss.n225 dvss.n130 6.61638
R805 dvss.n138 dvss.n137 6.48838
R806 dvss.n308 dvss.n307 6.25272
R807 dvss.n279 dvss.n278 6.24182
R808 dvss.n463 dvss.n454 5.62598
R809 dvss.n487 dvss.n478 5.62598
R810 dvss.n562 dvss.n561 5.62598
R811 dvss.n8 dvss.n2 5.62598
R812 dvss.n280 dvss.n279 5.45041
R813 dvss.n145 dvss.n144 5.36091
R814 dvss.n188 dvss.n154 5.32842
R815 dvss.n278 dvss.n276 5.14871
R816 dvss.n474 dvss.n473 4.81722
R817 dvss.n497 dvss.n496 4.81722
R818 dvss.n560 dvss.n14 4.81722
R819 dvss.n576 dvss.n575 4.81722
R820 dvss.n307 dvss.n306 4.13833
R821 dvss.n276 dvss.n275 3.91455
R822 dvss.n301 dvss.n76 3.78325
R823 dvss.n527 dvss.n526 3.6687
R824 dvss.n301 dvss.n300 3.64012
R825 dvss.n517 dvss.n39 3.4019
R826 dvss.n287 dvss.n286 3.38261
R827 dvss.n306 dvss.n68 3.20618
R828 dvss.n280 dvss.n77 2.68327
R829 dvss.n76 dvss.n75 2.51552
R830 dvss.n405 dvss.n335 2.25322
R831 dvss.n406 dvss.n405 2.25322
R832 dvss.n404 dvss.n402 2.25322
R833 dvss.n404 dvss.n403 2.25322
R834 dvss.n378 dvss.n377 2.25322
R835 dvss.n377 dvss.n357 2.25322
R836 dvss.n376 dvss.n362 2.25322
R837 dvss.n376 dvss.n375 2.25322
R838 dvss.n474 dvss.n453 2.25276
R839 dvss.n497 dvss.n477 2.25276
R840 dvss.n17 dvss.n14 2.25276
R841 dvss.n576 dvss.n1 2.25276
R842 dvss.n314 dvss.n313 2.11039
R843 dvss.n426 dvss.n421 1.86647
R844 dvss.n447 dvss.n446 1.70108
R845 dvss.n428 dvss.n427 1.60988
R846 dvss.n446 dvss.n445 1.59604
R847 dvss.n274 dvss.n55 1.58728
R848 dvss.t27 dvss.n532 1.50849
R849 dvss.n427 dvss.n426 1.38166
R850 dvss.n530 dvss.n529 1.30662
R851 dvss.n505 dvss.n504 1.23532
R852 dvss.n424 dvss.n422 1.2043
R853 dvss.n424 dvss.n423 1.2043
R854 dvss.n502 dvss.n0 1.08443
R855 dvss.n398 dvss.n335 1.03311
R856 dvss.n408 dvss.n406 1.03311
R857 dvss.n402 dvss.n401 1.03311
R858 dvss.n403 dvss.n333 1.03311
R859 dvss.n379 dvss.n378 1.03311
R860 dvss.n371 dvss.n357 1.03311
R861 dvss.n362 dvss.n361 1.03311
R862 dvss.n375 dvss.n374 1.03311
R863 dvss.n503 dvss.n502 0.979071
R864 dvss.n504 dvss.n503 0.978625
R865 dvss.n295 dvss.n294 0.878931
R866 dvss.n317 dvss.n316 0.780399
R867 dvss.n435 dvss.n434 0.7505
R868 dvss.n431 dvss.n430 0.714563
R869 dvss.n360 dvss.n359 0.709739
R870 dvss.n399 dvss.n397 0.709739
R871 dvss.n409 dvss.n332 0.709739
R872 dvss.n438 dvss.n437 0.688
R873 dvss.n429 dvss.n318 0.654856
R874 dvss.n44 dvss.n39 0.653561
R875 dvss.n358 dvss.n353 0.6255
R876 dvss.n380 dvss.n379 0.6255
R877 dvss.n351 dvss.n349 0.6255
R878 dvss.n384 dvss.n383 0.6255
R879 dvss.n347 dvss.n345 0.6255
R880 dvss.n388 dvss.n387 0.6255
R881 dvss.n343 dvss.n340 0.6255
R882 dvss.n392 dvss.n391 0.6255
R883 dvss.n396 dvss.n395 0.6255
R884 dvss.n401 dvss.n337 0.6255
R885 dvss.n333 dvss.n331 0.6255
R886 dvss.n412 dvss.n411 0.6255
R887 dvss.n329 dvss.n327 0.6255
R888 dvss.n416 dvss.n415 0.6255
R889 dvss.n365 dvss.n325 0.6255
R890 dvss.n368 dvss.n367 0.6255
R891 dvss.n371 dvss.n370 0.6255
R892 dvss.n439 dvss.n438 0.589954
R893 dvss.n431 dvss.n419 0.568435
R894 dvss.n507 dvss.n506 0.563319
R895 dvss.n146 dvss.n145 0.552784
R896 dvss.n224 dvss.n152 0.552784
R897 dvss.n150 dvss.n131 0.552784
R898 dvss.n154 dvss.n153 0.552784
R899 dvss.n430 dvss.n429 0.539326
R900 dvss.n440 dvss.n25 0.517167
R901 dvss.n433 dvss.n432 0.503217
R902 dvss.n434 dvss.n433 0.503217
R903 dvss.n436 dvss.n435 0.503217
R904 dvss.n437 dvss.n436 0.503217
R905 dvss.n426 dvss.n425 0.479667
R906 dvss.n427 dvss.n420 0.479667
R907 dvss.n452 dvss 0.472936
R908 dvss.n439 dvss.n318 0.466883
R909 dvss.n423 dvss.n421 0.451542
R910 dvss.n425 dvss.n424 0.451542
R911 dvss.n422 dvss.n420 0.451542
R912 dvss.n327 dvss.n326 0.440717
R913 dvss.n326 dvss.n325 0.440717
R914 dvss.n383 dvss.n350 0.440717
R915 dvss.n380 dvss.n350 0.440717
R916 dvss.n352 dvss.n351 0.440717
R917 dvss.n353 dvss.n352 0.440717
R918 dvss.n387 dvss.n346 0.440717
R919 dvss.n384 dvss.n346 0.440717
R920 dvss.n348 dvss.n347 0.440717
R921 dvss.n349 dvss.n348 0.440717
R922 dvss.n391 dvss.n342 0.440717
R923 dvss.n388 dvss.n342 0.440717
R924 dvss.n344 dvss.n343 0.440717
R925 dvss.n345 dvss.n344 0.440717
R926 dvss.n341 dvss.n337 0.440717
R927 dvss.n392 dvss.n341 0.440717
R928 dvss.n395 dvss.n339 0.440717
R929 dvss.n340 dvss.n339 0.440717
R930 dvss.n412 dvss.n328 0.440717
R931 dvss.n415 dvss.n328 0.440717
R932 dvss.n331 dvss.n330 0.440717
R933 dvss.n330 dvss.n329 0.440717
R934 dvss.n416 dvss.n324 0.440717
R935 dvss.n419 dvss.n324 0.440717
R936 dvss.n366 dvss.n365 0.440717
R937 dvss.n367 dvss.n366 0.440717
R938 dvss.n369 dvss.n368 0.440717
R939 dvss.n370 dvss.n369 0.440717
R940 dvss.n443 dvss.n442 0.40902
R941 dvss.n448 dvss.n443 0.40902
R942 dvss.n28 dvss.n26 0.38259
R943 dvss.n473 dvss.n454 0.379594
R944 dvss.n496 dvss.n478 0.379594
R945 dvss.n561 dvss.n560 0.379594
R946 dvss.n575 dvss.n2 0.379594
R947 dvss.n451 dvss.n450 0.377433
R948 dvss.n450 dvss.n449 0.377433
R949 dvss.n519 dvss.n515 0.366214
R950 dvss.n359 dvss.n358 0.359196
R951 dvss.n379 dvss.n354 0.359196
R952 dvss.n361 dvss.n354 0.359196
R953 dvss.n397 dvss.n396 0.359196
R954 dvss.n411 dvss.n332 0.359196
R955 dvss.n406 dvss.n334 0.359196
R956 dvss.n403 dvss.n334 0.359196
R957 dvss.n336 dvss.n335 0.359196
R958 dvss.n402 dvss.n336 0.359196
R959 dvss.n398 dvss.n338 0.359196
R960 dvss.n401 dvss.n338 0.359196
R961 dvss.n408 dvss.n407 0.359196
R962 dvss.n407 dvss.n333 0.359196
R963 dvss.n371 dvss.n364 0.359196
R964 dvss.n374 dvss.n364 0.359196
R965 dvss.n363 dvss.n357 0.359196
R966 dvss.n375 dvss.n363 0.359196
R967 dvss.n378 dvss.n356 0.359196
R968 dvss.n362 dvss.n356 0.359196
R969 dvss.n381 dvss.n353 0.351043
R970 dvss.n381 dvss.n380 0.351043
R971 dvss.n382 dvss.n351 0.351043
R972 dvss.n383 dvss.n382 0.351043
R973 dvss.n385 dvss.n349 0.351043
R974 dvss.n385 dvss.n384 0.351043
R975 dvss.n386 dvss.n347 0.351043
R976 dvss.n387 dvss.n386 0.351043
R977 dvss.n389 dvss.n345 0.351043
R978 dvss.n389 dvss.n388 0.351043
R979 dvss.n390 dvss.n343 0.351043
R980 dvss.n391 dvss.n390 0.351043
R981 dvss.n393 dvss.n340 0.351043
R982 dvss.n393 dvss.n392 0.351043
R983 dvss.n395 dvss.n394 0.351043
R984 dvss.n394 dvss.n337 0.351043
R985 dvss.n399 dvss.n398 0.351043
R986 dvss.n409 dvss.n408 0.351043
R987 dvss.n400 dvss.n396 0.351043
R988 dvss.n401 dvss.n400 0.351043
R989 dvss.n410 dvss.n333 0.351043
R990 dvss.n411 dvss.n410 0.351043
R991 dvss.n413 dvss.n331 0.351043
R992 dvss.n413 dvss.n412 0.351043
R993 dvss.n414 dvss.n329 0.351043
R994 dvss.n415 dvss.n414 0.351043
R995 dvss.n417 dvss.n327 0.351043
R996 dvss.n417 dvss.n416 0.351043
R997 dvss.n418 dvss.n325 0.351043
R998 dvss.n419 dvss.n418 0.351043
R999 dvss.n365 dvss.n323 0.351043
R1000 dvss.n367 dvss.n322 0.351043
R1001 dvss.n368 dvss.n321 0.351043
R1002 dvss.n370 dvss.n320 0.351043
R1003 dvss.n358 dvss.n355 0.351043
R1004 dvss.n379 dvss.n355 0.351043
R1005 dvss.n372 dvss.n371 0.351043
R1006 dvss.n361 dvss.n360 0.351043
R1007 dvss.n374 dvss.n373 0.351043
R1008 dvss.n475 dvss.n474 0.332643
R1009 dvss.n498 dvss.n497 0.332643
R1010 dvss.n500 dvss.n14 0.332643
R1011 dvss.n577 dvss.n576 0.332643
R1012 dvss.n441 dvss.n439 0.292684
R1013 dvss.n432 dvss.n323 0.288543
R1014 dvss.n434 dvss.n322 0.288543
R1015 dvss.n435 dvss.n321 0.288543
R1016 dvss.n437 dvss.n320 0.288543
R1017 dvss.n372 dvss.n319 0.288543
R1018 dvss.n373 dvss.n319 0.288543
R1019 dvss.n506 dvss.n505 0.2505
R1020 dvss.n475 dvss 0.242464
R1021 dvss.n498 dvss 0.242464
R1022 dvss.n500 dvss 0.242464
R1023 dvss dvss.n577 0.242464
R1024 dvss.n476 dvss.n475 0.224161
R1025 dvss.n499 dvss.n498 0.224161
R1026 dvss.n501 dvss.n500 0.224161
R1027 dvss.n577 dvss.n0 0.224161
R1028 dvss.n313 dvss.n56 0.217883
R1029 dvss.n441 dvss.n440 0.179826
R1030 dvss.n430 dvss.n428 0.1755
R1031 dvss.n432 dvss.n431 0.120065
R1032 dvss.n440 dvss 0.108642
R1033 dvss.n504 dvss.n476 0.106137
R1034 dvss.n503 dvss.n499 0.106137
R1035 dvss.n502 dvss.n501 0.106137
R1036 dvss.n452 dvss 0.038087
R1037 dvss.n508 dvss.n507 0.0357273
R1038 dvss.n507 dvss.n441 0.0153492
R1039 dvss.n505 dvss 0.0142289
R1040 dvss.n438 dvss.n319 0.00857584
R1041 dvss.n506 dvss.n452 0.000674014
R1042 multiplexer_0.vtrip_1.n0 multiplexer_0.vtrip_1.t0 41.2565
R1043 multiplexer_0.vtrip_1.n1 multiplexer_0.vtrip_1.n0 5.29988
R1044 multiplexer_0.vtrip_1.n1 multiplexer_0.vtrip_1.t12 16.8956
R1045 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.n11 17.2675
R1046 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.n1 1.62926
R1047 multiplexer_0.vtrip_1.n2 multiplexer_0.vtrip_1.n10 2.85792
R1048 multiplexer_0.vtrip_1.n4 multiplexer_0.vtrip_1.n2 3.14503
R1049 multiplexer_0.vtrip_1.n11 multiplexer_0.vtrip_1.n4 2.17823
R1050 multiplexer_0.vtrip_1.n11 multiplexer_0.vtrip_1.n6 0.967297
R1051 multiplexer_0.vtrip_1.n6 multiplexer_0.vtrip_1.n8 2.84816
R1052 multiplexer_0.vtrip_1.n10 multiplexer_0.vtrip_1.t4 97.2843
R1053 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.n9 0.171398
R1054 multiplexer_0.vtrip_1.n10 multiplexer_0.vtrip_1.n9 0.162609
R1055 multiplexer_0.vtrip_1.n9 multiplexer_0.vtrip_1 3.32193
R1056 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.t6 18.1873
R1057 multiplexer_0.vtrip_1.n8 multiplexer_0.vtrip_1.t11 97.2843
R1058 multiplexer_0.vtrip_1.n8 multiplexer_0.vtrip_1 3.4938
R1059 multiplexer_0.vtrip_1.t8 multiplexer_0.vtrip_1 18.5516
R1060 multiplexer_0.vtrip_1.n6 multiplexer_0.vtrip_1 3.32193
R1061 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.n7 1.67907
R1062 multiplexer_0.vtrip_1.t9 multiplexer_0.vtrip_1.n7 16.8731
R1063 multiplexer_0.vtrip_1.n7 multiplexer_0.vtrip_1.t2 16.5088
R1064 multiplexer_0.vtrip_1.n4 multiplexer_0.vtrip_1 3.32193
R1065 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.n5 1.67907
R1066 multiplexer_0.vtrip_1.t3 multiplexer_0.vtrip_1.n5 16.8731
R1067 multiplexer_0.vtrip_1.n5 multiplexer_0.vtrip_1.t5 16.5088
R1068 multiplexer_0.vtrip_1.n2 multiplexer_0.vtrip_1 3.32193
R1069 multiplexer_0.vtrip_1 multiplexer_0.vtrip_1.n3 1.67907
R1070 multiplexer_0.vtrip_1.t7 multiplexer_0.vtrip_1.n3 16.8731
R1071 multiplexer_0.vtrip_1.n3 multiplexer_0.vtrip_1.t10 16.5088
R1072 multiplexer_0.vtrip_1.n0 multiplexer_0.vtrip_1.t1 227.385
R1073 multiplexer_0.trans_gate_m_29.in.t1 multiplexer_0.trans_gate_m_29.in.n0 228.216
R1074 multiplexer_0.trans_gate_m_29.in.n5 multiplexer_0.trans_gate_m_29.in.n0 1.5005
R1075 multiplexer_0.trans_gate_m_29.in.n0 multiplexer_0.trans_gate_m_29.in.t0 83.695
R1076 multiplexer_0.trans_gate_m_29.in multiplexer_0.trans_gate_m_29.in.n5 0.104667
R1077 multiplexer_0.trans_gate_m_29.in.n5 multiplexer_0.trans_gate_m_29.in.n4 4.43682
R1078 multiplexer_0.trans_gate_m_29.in.n2 multiplexer_0.trans_gate_m_29.in.n1 1.5005
R1079 multiplexer_0.trans_gate_m_29.in multiplexer_0.trans_gate_m_29.in.n2 0.104667
R1080 multiplexer_0.trans_gate_m_29.in.n4 multiplexer_0.trans_gate_m_29.in.n2 0.459875
R1081 multiplexer_0.trans_gate_m_29.in.n4 multiplexer_0.trans_gate_m_29.in 0.564042
R1082 multiplexer_0.trans_gate_m_29.in multiplexer_0.trans_gate_m_29.in.n3 1.60467
R1083 multiplexer_0.trans_gate_m_29.in.n3 multiplexer_0.trans_gate_m_29.in.t5 83.695
R1084 multiplexer_0.trans_gate_m_29.in.n3 multiplexer_0.trans_gate_m_29.in.t3 228.216
R1085 multiplexer_0.trans_gate_m_29.in.n1 multiplexer_0.trans_gate_m_29.in.t2 83.695
R1086 multiplexer_0.trans_gate_m_29.in.n1 multiplexer_0.trans_gate_m_29.in.t4 228.216
R1087 multiplexer_0.trans_gate_m_31.out.t1 multiplexer_0.trans_gate_m_31.out.n0 228.216
R1088 multiplexer_0.trans_gate_m_31.out.n5 multiplexer_0.trans_gate_m_31.out.n0 1.5005
R1089 multiplexer_0.trans_gate_m_31.out.n0 multiplexer_0.trans_gate_m_31.out.t4 83.695
R1090 multiplexer_0.trans_gate_m_31.out multiplexer_0.trans_gate_m_31.out.n5 0.104667
R1091 multiplexer_0.trans_gate_m_31.out.n5 multiplexer_0.trans_gate_m_31.out.n3 0.459875
R1092 multiplexer_0.trans_gate_m_31.out.n3 multiplexer_0.trans_gate_m_31.out 0.553625
R1093 multiplexer_0.trans_gate_m_31.out multiplexer_0.trans_gate_m_31.out.n4 1.60467
R1094 multiplexer_0.trans_gate_m_31.out.n4 multiplexer_0.trans_gate_m_31.out.t0 83.695
R1095 multiplexer_0.trans_gate_m_31.out.n4 multiplexer_0.trans_gate_m_31.out.t5 228.216
R1096 multiplexer_0.trans_gate_m_31.out.n3 multiplexer_0.trans_gate_m_31.out.n2 4.43682
R1097 multiplexer_0.trans_gate_m_31.out.n2 multiplexer_0.trans_gate_m_31.out.n1 1.5005
R1098 multiplexer_0.trans_gate_m_31.out multiplexer_0.trans_gate_m_31.out.n2 0.104667
R1099 multiplexer_0.trans_gate_m_31.out.n1 multiplexer_0.trans_gate_m_31.out.t2 83.695
R1100 multiplexer_0.trans_gate_m_31.out.n1 multiplexer_0.trans_gate_m_31.out.t3 228.216
R1101 avss.n734 avss.n113 52837.8
R1102 avss.n734 avss.n114 52837.8
R1103 avss.n735 avss.n114 52837.8
R1104 avss.n735 avss.n113 52837.8
R1105 avss.n485 avss.n137 10442.2
R1106 avss.n612 avss.n249 6744.4
R1107 avss.n418 avss.n253 6744.4
R1108 avss.n612 avss.n253 6744.4
R1109 avss.n377 avss.n356 6744.4
R1110 avss.n418 avss.n377 6744.4
R1111 avss.n571 avss.n356 6744.4
R1112 avss.n571 avss.n317 6744.4
R1113 avss.n636 avss.n635 6328.99
R1114 avss.n487 avss.n214 6328.99
R1115 avss.n636 avss.n214 6328.99
R1116 avss.n647 avss.n168 6227.45
R1117 avss.n272 avss.n239 6216.37
R1118 avss.n623 avss.n235 6216.37
R1119 avss.n623 avss.n239 6216.37
R1120 avss.n557 avss.n429 6216.37
R1121 avss.n429 avss.n235 6216.37
R1122 avss.n557 avss.n431 6216.37
R1123 avss.n489 avss.n431 6216.37
R1124 avss.n656 avss.n137 6184.38
R1125 avss.n488 avss.n486 4558.19
R1126 avss.n485 avss.n484 3690.48
R1127 avss.n488 avss.n487 3618.39
R1128 avss.n657 avss.n656 3386.05
R1129 avss.n489 avss.n488 3228.89
R1130 avss.n729 avss.n118 3052.71
R1131 avss.n728 avss.n118 3052.71
R1132 avss.n728 avss.n117 3052.71
R1133 avss.n729 avss.n117 3052.71
R1134 avss.n162 avss.n137 2992.39
R1135 avss.n158 avss.n157 2723.4
R1136 avss.n157 avss.n134 2723.4
R1137 avss.n712 avss.n141 2723.4
R1138 avss.n693 avss.n141 2723.4
R1139 avss.n153 avss.n151 2723.4
R1140 avss.n151 avss.n135 2723.4
R1141 avss.n154 avss.n140 2723.4
R1142 avss.n695 avss.n154 2723.4
R1143 avss.n674 avss.n159 2723.4
R1144 avss.n674 avss.n136 2723.4
R1145 avss.n669 avss.n139 2723.4
R1146 avss.n687 avss.n669 2723.4
R1147 avss.n160 avss.n133 2723.4
R1148 avss.n714 avss.n133 2723.4
R1149 avss.n659 avss.n138 2723.4
R1150 avss.n668 avss.n659 2723.4
R1151 avss.n486 avss.n485 2564.43
R1152 avss.t217 avss.n502 2496.57
R1153 avss.t217 avss.n503 2496.57
R1154 avss.n430 avss.t148 2496.57
R1155 avss.n570 avss.t148 2496.57
R1156 avss.t157 avss.n572 2496.57
R1157 avss.t157 avss.n318 2496.57
R1158 avss.n483 avss.t246 2496.57
R1159 avss.n476 avss.t246 2496.57
R1160 avss.n195 avss.t254 2496.57
R1161 avss.n201 avss.t254 2496.57
R1162 avss.t216 avss.n544 2496.57
R1163 avss.t216 avss.n545 2496.57
R1164 avss.n428 avss.t136 2496.57
R1165 avss.n376 avss.t136 2496.57
R1166 avss.t191 avss.n398 2496.57
R1167 avss.t191 avss.n319 2496.57
R1168 avss.t214 avss.n234 2496.57
R1169 avss.t214 avss.n624 2496.57
R1170 avss.n622 avss.t101 2496.57
R1171 avss.n252 avss.t101 2496.57
R1172 avss.t30 avss.n408 2496.57
R1173 avss.t30 avss.n320 2496.57
R1174 avss.n633 avss.t187 2496.57
R1175 avss.n238 avss.t187 2496.57
R1176 avss.t197 avss.n248 2496.57
R1177 avss.t197 avss.n613 2496.57
R1178 avss.n611 avss.t151 2496.57
R1179 avss.n323 avss.t151 2496.57
R1180 avss.t112 avss.n513 2496.57
R1181 avss.t112 avss.n514 2496.57
R1182 avss.t239 avss.n373 2496.57
R1183 avss.t239 avss.n419 2496.57
R1184 avss.n417 avss.t47 2496.57
R1185 avss.t47 avss.n324 2496.57
R1186 avss.n500 avss.t188 2496.57
R1187 avss.n556 avss.t188 2496.57
R1188 avss.t182 avss.n558 2496.57
R1189 avss.t182 avss.n559 2496.57
R1190 avss.t29 avss.n388 2496.57
R1191 avss.t29 avss.n325 2496.57
R1192 avss.t186 avss.n440 2496.57
R1193 avss.t186 avss.n490 2496.57
R1194 avss.t57 avss.n441 2496.57
R1195 avss.t57 avss.n450 2496.57
R1196 avss.n329 avss.t196 2496.57
R1197 avss.n583 avss.t196 2496.57
R1198 avss.n582 avss.n326 2394.09
R1199 avss.n582 avss.n327 2394.09
R1200 avss.n330 avss.n327 2394.09
R1201 avss.n330 avss.n326 2394.09
R1202 avss.n451 avss.n449 2394.09
R1203 avss.n452 avss.n449 2394.09
R1204 avss.n452 avss.n447 2394.09
R1205 avss.n451 avss.n447 2394.09
R1206 avss.n491 avss.n439 2394.09
R1207 avss.n492 avss.n439 2394.09
R1208 avss.n492 avss.n437 2394.09
R1209 avss.n491 avss.n437 2394.09
R1210 avss.n389 avss.n387 2394.09
R1211 avss.n390 avss.n387 2394.09
R1212 avss.n390 avss.n385 2394.09
R1213 avss.n389 avss.n385 2394.09
R1214 avss.n560 avss.n364 2394.09
R1215 avss.n561 avss.n364 2394.09
R1216 avss.n561 avss.n362 2394.09
R1217 avss.n560 avss.n362 2394.09
R1218 avss.n555 avss.n432 2394.09
R1219 avss.n555 avss.n433 2394.09
R1220 avss.n435 avss.n433 2394.09
R1221 avss.n435 avss.n432 2394.09
R1222 avss.n381 avss.n378 2394.09
R1223 avss.n381 avss.n379 2394.09
R1224 avss.n416 avss.n379 2394.09
R1225 avss.n416 avss.n378 2394.09
R1226 avss.n420 avss.n372 2394.09
R1227 avss.n421 avss.n372 2394.09
R1228 avss.n421 avss.n370 2394.09
R1229 avss.n420 avss.n370 2394.09
R1230 avss.n515 avss.n512 2394.09
R1231 avss.n516 avss.n512 2394.09
R1232 avss.n516 avss.n510 2394.09
R1233 avss.n515 avss.n510 2394.09
R1234 avss.n322 avss.n254 2394.09
R1235 avss.n322 avss.n255 2394.09
R1236 avss.n610 avss.n255 2394.09
R1237 avss.n610 avss.n254 2394.09
R1238 avss.n614 avss.n247 2394.09
R1239 avss.n615 avss.n247 2394.09
R1240 avss.n615 avss.n245 2394.09
R1241 avss.n614 avss.n245 2394.09
R1242 avss.n237 avss.n226 2394.09
R1243 avss.n237 avss.n227 2394.09
R1244 avss.n632 avss.n227 2394.09
R1245 avss.n632 avss.n226 2394.09
R1246 avss.n596 avss.n316 2394.09
R1247 avss.n595 avss.n316 2394.09
R1248 avss.n595 avss.n259 2394.09
R1249 avss.n596 avss.n259 2394.09
R1250 avss.n308 avss.n269 2394.09
R1251 avss.n308 avss.n270 2394.09
R1252 avss.n303 avss.n270 2394.09
R1253 avss.n303 avss.n269 2394.09
R1254 avss.n287 avss.n280 2394.09
R1255 avss.n287 avss.n281 2394.09
R1256 avss.n283 avss.n281 2394.09
R1257 avss.n283 avss.n280 2394.09
R1258 avss.n409 avss.n407 2394.09
R1259 avss.n410 avss.n407 2394.09
R1260 avss.n410 avss.n405 2394.09
R1261 avss.n409 avss.n405 2394.09
R1262 avss.n251 avss.n240 2394.09
R1263 avss.n251 avss.n241 2394.09
R1264 avss.n621 avss.n241 2394.09
R1265 avss.n621 avss.n240 2394.09
R1266 avss.n625 avss.n233 2394.09
R1267 avss.n626 avss.n233 2394.09
R1268 avss.n626 avss.n231 2394.09
R1269 avss.n625 avss.n231 2394.09
R1270 avss.n399 avss.n397 2394.09
R1271 avss.n400 avss.n397 2394.09
R1272 avss.n400 avss.n395 2394.09
R1273 avss.n399 avss.n395 2394.09
R1274 avss.n375 avss.n365 2394.09
R1275 avss.n375 avss.n366 2394.09
R1276 avss.n427 avss.n366 2394.09
R1277 avss.n427 avss.n365 2394.09
R1278 avss.n546 avss.n524 2394.09
R1279 avss.n547 avss.n524 2394.09
R1280 avss.n547 avss.n522 2394.09
R1281 avss.n546 avss.n522 2394.09
R1282 avss.n200 avss.n192 2394.09
R1283 avss.n200 avss.n193 2394.09
R1284 avss.n196 avss.n193 2394.09
R1285 avss.n196 avss.n192 2394.09
R1286 avss.n477 avss.n473 2394.09
R1287 avss.n477 avss.n474 2394.09
R1288 avss.n482 avss.n474 2394.09
R1289 avss.n482 avss.n473 2394.09
R1290 avss.n573 avss.n355 2394.09
R1291 avss.n574 avss.n355 2394.09
R1292 avss.n574 avss.n353 2394.09
R1293 avss.n573 avss.n353 2394.09
R1294 avss.n569 avss.n357 2394.09
R1295 avss.n569 avss.n358 2394.09
R1296 avss.n360 avss.n358 2394.09
R1297 avss.n360 avss.n357 2394.09
R1298 avss.n504 avss.n499 2394.09
R1299 avss.n505 avss.n499 2394.09
R1300 avss.n505 avss.n497 2394.09
R1301 avss.n504 avss.n497 2394.09
R1302 avss.n212 avss.n203 2394.09
R1303 avss.n212 avss.n204 2394.09
R1304 avss.n207 avss.n204 2394.09
R1305 avss.n207 avss.n203 2394.09
R1306 avss.n649 avss.n163 2394.09
R1307 avss.n649 avss.n164 2394.09
R1308 avss.n653 avss.n164 2394.09
R1309 avss.n653 avss.n163 2394.09
R1310 avss.n223 avss.n216 2394.09
R1311 avss.n223 avss.n217 2394.09
R1312 avss.n219 avss.n217 2394.09
R1313 avss.n219 avss.n216 2394.09
R1314 avss.n190 avss.n188 2394.09
R1315 avss.n638 avss.n190 2394.09
R1316 avss.n639 avss.n638 2394.09
R1317 avss.n639 avss.n188 2394.09
R1318 avss.n503 avss.n431 2027.45
R1319 avss.n431 avss.n430 2027.45
R1320 avss.n545 avss.n429 2027.45
R1321 avss.n429 avss.n428 2027.45
R1322 avss.n624 avss.n623 2027.45
R1323 avss.n623 avss.n622 2027.45
R1324 avss.n239 avss.n238 2027.45
R1325 avss.n248 avss.n239 2027.45
R1326 avss.n514 avss.n235 2027.45
R1327 avss.n373 avss.n235 2027.45
R1328 avss.n557 avss.n556 2027.45
R1329 avss.n558 avss.n557 2027.45
R1330 avss.n490 avss.n489 2027.45
R1331 avss.n489 avss.n441 2027.45
R1332 avss.n484 avss.n162 2007.05
R1333 avss.n655 avss.n162 1963.94
R1334 avss.n571 avss.n570 1908.82
R1335 avss.n572 avss.n571 1908.82
R1336 avss.n377 avss.n376 1908.82
R1337 avss.n398 avss.n377 1908.82
R1338 avss.n253 avss.n252 1908.82
R1339 avss.n408 avss.n253 1908.82
R1340 avss.n613 avss.n612 1908.82
R1341 avss.n612 avss.n611 1908.82
R1342 avss.n419 avss.n418 1908.82
R1343 avss.n418 avss.n417 1908.82
R1344 avss.n559 avss.n356 1908.82
R1345 avss.n388 avss.n356 1908.82
R1346 avss.n450 avss.n317 1908.82
R1347 avss.n329 avss.n317 1908.82
R1348 avss.n489 avss.n317 1784.13
R1349 avss.n311 avss.n263 1552.82
R1350 avss.n603 avss.n263 1552.82
R1351 avss.n600 avss.n265 1552.82
R1352 avss.n601 avss.n600 1552.82
R1353 avss.n295 avss.n279 1552.82
R1354 avss.n295 avss.n273 1552.82
R1355 avss.n292 avss.n274 1552.82
R1356 avss.n300 avss.n274 1552.82
R1357 avss.n341 avss.n338 1552.82
R1358 avss.n338 avss.n337 1552.82
R1359 avss.n347 avss.n343 1552.82
R1360 avss.n347 avss.n344 1552.82
R1361 avss.n462 avss.n459 1552.82
R1362 avss.n459 avss.n442 1552.82
R1363 avss.n465 avss.n443 1552.82
R1364 avss.n471 avss.n443 1552.82
R1365 avss.n542 avss.n525 1552.82
R1366 avss.n531 avss.n525 1552.82
R1367 avss.n536 avss.n191 1552.82
R1368 avss.n646 avss.n173 1552.82
R1369 avss.n646 avss.n174 1552.82
R1370 avss.n181 avss.n166 1552.82
R1371 avss.n590 avss.n584 1552.82
R1372 avss.n586 avss.n584 1552.82
R1373 avss.n587 avss.n586 1552.82
R1374 avss.n590 avss.n587 1552.82
R1375 avss.n689 avss.n688 1524.71
R1376 avss.n688 avss.n142 1524.71
R1377 avss.n698 avss.n696 1524.71
R1378 avss.n698 avss.n697 1524.71
R1379 avss.n683 avss.n670 1524.71
R1380 avss.n683 avss.n682 1524.71
R1381 avss.n664 avss.n660 1524.71
R1382 avss.n664 avss.n132 1524.71
R1383 avss.n592 avss.n317 1481.39
R1384 avss.n476 avss.n169 1380.39
R1385 avss.n202 avss.n201 1380.39
R1386 avss.n733 avss.n112 1306.82
R1387 avss.n733 avss.n732 1306.74
R1388 avss.n195 avss.n170 1267.16
R1389 avss.n487 avss.n440 1266.54
R1390 avss.n655 avss.n161 1248.77
R1391 avss.n544 avss.n543 1218.63
R1392 avss.n689 avss.n158 1198.69
R1393 avss.n712 avss.n142 1198.69
R1394 avss.n142 avss.n134 1198.69
R1395 avss.n693 avss.n689 1198.69
R1396 avss.n696 avss.n153 1198.69
R1397 avss.n697 avss.n140 1198.69
R1398 avss.n697 avss.n135 1198.69
R1399 avss.n696 avss.n695 1198.69
R1400 avss.n670 avss.n159 1198.69
R1401 avss.n682 avss.n139 1198.69
R1402 avss.n682 avss.n136 1198.69
R1403 avss.n687 avss.n670 1198.69
R1404 avss.n660 avss.n160 1198.69
R1405 avss.n138 avss.n132 1198.69
R1406 avss.n714 avss.n132 1198.69
R1407 avss.n668 avss.n660 1198.69
R1408 avss.n656 avss.n655 1183.26
R1409 avss.n647 avss.n166 957.487
R1410 avss.n636 avss.n191 929.78
R1411 avss.n486 avss.n168 881.452
R1412 avss.t25 avss.n167 839.736
R1413 avss.t25 avss.n637 839.736
R1414 avss.n206 avss.t26 839.736
R1415 avss.n213 avss.t26 839.736
R1416 avss.n736 avss.n112 815.148
R1417 avss.n311 avss.n268 799.588
R1418 avss.n268 avss.n265 799.588
R1419 avss.n601 avss.n262 799.588
R1420 avss.n603 avss.n262 799.588
R1421 avss.n293 avss.n279 799.588
R1422 avss.n293 avss.n292 799.588
R1423 avss.n300 avss.n275 799.588
R1424 avss.n275 avss.n273 799.588
R1425 avss.n341 avss.n334 799.588
R1426 avss.n343 avss.n334 799.588
R1427 avss.n344 avss.n335 799.588
R1428 avss.n337 avss.n335 799.588
R1429 avss.n466 avss.n462 799.588
R1430 avss.n466 avss.n465 799.588
R1431 avss.n471 avss.n444 799.588
R1432 avss.n444 avss.n442 799.588
R1433 avss.n542 avss.n526 799.588
R1434 avss.n531 avss.n530 799.588
R1435 avss.n530 avss.n191 799.588
R1436 avss.n538 avss.n526 799.588
R1437 avss.n173 avss.n172 799.588
R1438 avss.n180 avss.n174 799.588
R1439 avss.n183 avss.n180 799.588
R1440 avss.n172 avss.n166 799.588
R1441 avss.n268 avss.n267 753.236
R1442 avss.n267 avss.n262 753.236
R1443 avss.n294 avss.n293 753.236
R1444 avss.n294 avss.n275 753.236
R1445 avss.n348 avss.n334 753.236
R1446 avss.n348 avss.n335 753.236
R1447 avss.n467 avss.n466 753.236
R1448 avss.n467 avss.n444 753.236
R1449 avss.n530 avss.n529 753.236
R1450 avss.n529 avss.n526 753.236
R1451 avss.n172 avss.n171 753.236
R1452 avss.n180 avss.n171 753.236
R1453 avss.t147 avss.n336 720.404
R1454 avss.n464 avss.t189 720.404
R1455 avss.n489 avss.n472 709.321
R1456 avss.t161 avss.n170 700.981
R1457 avss.n543 avss.t141 700.981
R1458 avss.n206 avss.n168 680.133
R1459 avss.n637 avss.n636 672.878
R1460 avss.n214 avss.n213 672.878
R1461 avss.n732 avss.n731 663.183
R1462 avss.n647 avss.n169 647.059
R1463 avss.n654 avss.t41 632.672
R1464 avss.n648 avss.t41 632.672
R1465 avss.n636 avss.n202 620.098
R1466 avss.n342 avss.n317 609.572
R1467 avss.n647 avss.n167 554.909
R1468 avss.n538 avss.n537 550.293
R1469 avss.n183 avss.n182 550.293
R1470 avss.n648 avss.n647 513.789
R1471 avss.n502 avss.n501 512.255
R1472 avss.n592 avss.n318 512.255
R1473 avss.n484 avss.n483 512.255
R1474 avss.n592 avss.n319 512.255
R1475 avss.n234 avss.n215 512.255
R1476 avss.n592 avss.n320 512.255
R1477 avss.n634 avss.n633 512.255
R1478 avss.n592 avss.n323 512.255
R1479 avss.n513 avss.n215 512.255
R1480 avss.n592 avss.n324 512.255
R1481 avss.n501 avss.n500 512.255
R1482 avss.n592 avss.n325 512.255
R1483 avss.n592 avss.n583 512.255
R1484 avss.n636 avss.n215 500.577
R1485 avss.n501 avss.n214 500.577
R1486 avss.n658 avss.n657 447.11
R1487 avss.t215 avss.n225 426.997
R1488 avss.n288 avss.t215 426.997
R1489 avss.n302 avss.t158 426.997
R1490 avss.n309 avss.t158 426.997
R1491 avss.t61 avss.n264 426.997
R1492 avss.t61 avss.n593 426.997
R1493 avss.t13 avss 380.286
R1494 avss.t10 avss 380.286
R1495 avss.t5 avss 380.286
R1496 avss.t60 avss.n161 319.26
R1497 avss.n224 avss.t60 319.26
R1498 avss avss.t13 296.784
R1499 avss.t10 avss 296.784
R1500 avss avss.t5 296.784
R1501 avss.n349 avss.n348 292.5
R1502 avss.n348 avss.t147 292.5
R1503 avss.n344 avss.n331 292.5
R1504 avss.n344 avss.n336 292.5
R1505 avss.n337 avss.n332 292.5
R1506 avss.n337 avss.n336 292.5
R1507 avss.n339 avss.n338 292.5
R1508 avss.t147 avss.n338 292.5
R1509 avss.n341 avss.n340 292.5
R1510 avss.n342 avss.n341 292.5
R1511 avss.n345 avss.n343 292.5
R1512 avss.n343 avss.n342 292.5
R1513 avss.n347 avss.n346 292.5
R1514 avss.t147 avss.n347 292.5
R1515 avss.n468 avss.n467 292.5
R1516 avss.n467 avss.t189 292.5
R1517 avss.n471 avss.n470 292.5
R1518 avss.n472 avss.n471 292.5
R1519 avss.n457 avss.n442 292.5
R1520 avss.n472 avss.n442 292.5
R1521 avss.n460 avss.n459 292.5
R1522 avss.n459 avss.t189 292.5
R1523 avss.n462 avss.n461 292.5
R1524 avss.n464 avss.n462 292.5
R1525 avss.n465 avss.n463 292.5
R1526 avss.n465 avss.n464 292.5
R1527 avss.n445 avss.n443 292.5
R1528 avss.n443 avss.t189 292.5
R1529 avss.n539 avss.n538 292.5
R1530 avss.n536 avss.n535 292.5
R1531 avss.n534 avss.n191 292.5
R1532 avss.n178 avss.n166 292.5
R1533 avss.n181 avss.n179 292.5
R1534 avss.n184 avss.n183 292.5
R1535 avss.n176 avss.n171 292.5
R1536 avss.t161 avss.n171 292.5
R1537 avss.n644 avss.n174 292.5
R1538 avss.n174 avss.n170 292.5
R1539 avss.n175 avss.n173 292.5
R1540 avss.n173 avss.n169 292.5
R1541 avss.n646 avss.n645 292.5
R1542 avss.t161 avss.n646 292.5
R1543 avss.n529 avss.n528 292.5
R1544 avss.n529 avss.t141 292.5
R1545 avss.n542 avss.n541 292.5
R1546 avss.n543 avss.n542 292.5
R1547 avss.n532 avss.n531 292.5
R1548 avss.n531 avss.n202 292.5
R1549 avss.n527 avss.n525 292.5
R1550 avss.n525 avss.t141 292.5
R1551 avss.n294 avss.n277 292.5
R1552 avss.t44 avss.n294 292.5
R1553 avss.n300 avss.n299 292.5
R1554 avss.n301 avss.n300 292.5
R1555 avss.n297 avss.n273 292.5
R1556 avss.n301 avss.n273 292.5
R1557 avss.n296 avss.n295 292.5
R1558 avss.n295 avss.t44 292.5
R1559 avss.n279 avss.n278 292.5
R1560 avss.n289 avss.n279 292.5
R1561 avss.n292 avss.n291 292.5
R1562 avss.n292 avss.n289 292.5
R1563 avss.n276 avss.n274 292.5
R1564 avss.t44 avss.n274 292.5
R1565 avss.n267 avss.n260 292.5
R1566 avss.n267 avss.t73 292.5
R1567 avss.n601 avss.n258 292.5
R1568 avss.n602 avss.n601 292.5
R1569 avss.n604 avss.n603 292.5
R1570 avss.n603 avss.n602 292.5
R1571 avss.n266 avss.n263 292.5
R1572 avss.t73 avss.n263 292.5
R1573 avss.n312 avss.n311 292.5
R1574 avss.n311 avss.n310 292.5
R1575 avss.n314 avss.n265 292.5
R1576 avss.n310 avss.n265 292.5
R1577 avss.n600 avss.n599 292.5
R1578 avss.n600 avss.t73 292.5
R1579 avss.n590 avss.n589 292.5
R1580 avss.n591 avss.n590 292.5
R1581 avss.n588 avss.n584 292.5
R1582 avss.n584 avss.t152 292.5
R1583 avss.n586 avss.n123 292.5
R1584 avss.n586 avss.n585 292.5
R1585 avss.n587 avss.n122 292.5
R1586 avss.n587 avss.t152 292.5
R1587 avss.n581 avss.n328 278.212
R1588 avss.n354 avss.n352 278.212
R1589 avss.n386 avss.n384 278.212
R1590 avss.n396 avss.n394 278.212
R1591 avss.n382 avss.n380 278.212
R1592 avss.n406 avss.n404 278.212
R1593 avss.n321 avss.n256 278.212
R1594 avss.n597 avss.n315 278.212
R1595 avss.n448 avss.n446 278.212
R1596 avss.n568 avss.n359 278.212
R1597 avss.n363 avss.n361 278.212
R1598 avss.n374 avss.n367 278.212
R1599 avss.n371 avss.n369 278.212
R1600 avss.n250 avss.n242 278.212
R1601 avss.n246 avss.n244 278.212
R1602 avss.n307 avss.n271 278.212
R1603 avss.n478 avss.n475 278.212
R1604 avss.n650 avss.n165 278.212
R1605 avss.n438 avss.n436 278.212
R1606 avss.n498 avss.n496 278.212
R1607 avss.n554 avss.n434 278.212
R1608 avss.n523 avss.n521 278.212
R1609 avss.n511 avss.n509 278.212
R1610 avss.n232 avss.n230 278.212
R1611 avss.n236 avss.n228 278.212
R1612 avss.n286 avss.n282 278.212
R1613 avss.n222 avss.n218 278.212
R1614 avss.n211 avss.n205 278.212
R1615 avss.n199 avss.n194 278.212
R1616 avss.n189 avss.n186 278.212
R1617 avss.n635 avss.n224 255.822
R1618 avss.n713 avss.t31 241.147
R1619 avss.n302 avss.n301 228.715
R1620 avss.t14 avss 226.321
R1621 avss.n289 avss.n288 225.026
R1622 avss.n310 avss.n309 225.026
R1623 avss.n694 avss.n658 220.312
R1624 avss.n581 avss.n580 214.03
R1625 avss.n575 avss.n354 214.03
R1626 avss.n391 avss.n386 214.03
R1627 avss.n401 avss.n396 214.03
R1628 avss.n383 avss.n382 214.03
R1629 avss.n411 avss.n406 214.03
R1630 avss.n321 avss.n257 214.03
R1631 avss.n594 avss.n315 214.03
R1632 avss.n453 avss.n448 214.03
R1633 avss.n568 avss.n567 214.03
R1634 avss.n562 avss.n363 214.03
R1635 avss.n374 avss.n368 214.03
R1636 avss.n422 avss.n371 214.03
R1637 avss.n250 avss.n243 214.03
R1638 avss.n616 avss.n246 214.03
R1639 avss.n307 avss.n306 214.03
R1640 avss.n479 avss.n478 214.03
R1641 avss.n651 avss.n650 214.03
R1642 avss.n493 avss.n438 214.03
R1643 avss.n506 avss.n498 214.03
R1644 avss.n554 avss.n553 214.03
R1645 avss.n548 avss.n523 214.03
R1646 avss.n517 avss.n511 214.03
R1647 avss.n627 avss.n232 214.03
R1648 avss.n236 avss.n229 214.03
R1649 avss.n286 avss.n285 214.03
R1650 avss.n222 avss.n221 214.03
R1651 avss.n211 avss.n210 214.03
R1652 avss.n199 avss.n198 214.03
R1653 avss.n189 avss.n187 214.03
R1654 avss.n579 avss.n328 204.909
R1655 avss.n576 avss.n352 204.909
R1656 avss.n392 avss.n384 204.909
R1657 avss.n402 avss.n394 204.909
R1658 avss.n415 avss.n380 204.909
R1659 avss.n412 avss.n404 204.909
R1660 avss.n609 avss.n256 204.909
R1661 avss.n454 avss.n446 204.909
R1662 avss.n566 avss.n359 204.909
R1663 avss.n563 avss.n361 204.909
R1664 avss.n426 avss.n367 204.909
R1665 avss.n423 avss.n369 204.909
R1666 avss.n620 avss.n242 204.909
R1667 avss.n617 avss.n244 204.909
R1668 avss.n305 avss.n271 204.909
R1669 avss.n481 avss.n475 204.909
R1670 avss.n652 avss.n165 204.909
R1671 avss.n494 avss.n436 204.909
R1672 avss.n507 avss.n496 204.909
R1673 avss.n552 avss.n434 204.909
R1674 avss.n549 avss.n521 204.909
R1675 avss.n518 avss.n509 204.909
R1676 avss.n628 avss.n230 204.909
R1677 avss.n631 avss.n228 204.909
R1678 avss.n284 avss.n282 204.909
R1679 avss.n220 avss.n218 204.909
R1680 avss.n209 avss.n205 204.909
R1681 avss.n197 avss.n194 204.909
R1682 avss.n640 avss.n186 204.909
R1683 avss.n635 avss.n634 190.315
R1684 avss.n602 avss.n264 188.137
R1685 avss.n598 avss.n597 187.107
R1686 avss.n655 avss.n654 183.107
R1687 avss.n691 avss.n144 174.306
R1688 avss.n710 avss.n144 174.306
R1689 avss.n699 avss.n150 174.306
R1690 avss.n700 avss.n699 174.306
R1691 avss.n685 avss.n684 174.306
R1692 avss.n684 avss.n681 174.306
R1693 avss.n666 avss.n665 174.306
R1694 avss.n665 avss.n131 174.306
R1695 avss.n711 avss.n143 170.748
R1696 avss.n692 avss.n143 170.748
R1697 avss.n155 avss.n149 170.748
R1698 avss.n156 avss.n155 170.748
R1699 avss.n673 avss.n671 170.748
R1700 avss.n686 avss.n671 170.748
R1701 avss.n662 avss.n661 170.748
R1702 avss.n667 avss.n662 170.748
R1703 avss.n690 avss.n145 166.988
R1704 avss.n152 avss.n148 166.988
R1705 avss.n675 avss.n672 166.988
R1706 avss.n663 avss.n130 166.988
R1707 avss.n709 avss.n708 166.934
R1708 avss.n702 avss.n701 166.934
R1709 avss.n680 avss.n679 166.934
R1710 avss.n716 avss.n715 166.934
R1711 avss.n537 avss.n536 158.911
R1712 avss.n182 avss.n181 158.911
R1713 avss.t0 avss.n114 145.641
R1714 avss.n120 avss.t14 143.45
R1715 avss avss.t0 142.819
R1716 avss.n711 avss.n710 141.554
R1717 avss.n692 avss.n691 141.554
R1718 avss.n691 avss.n690 141.554
R1719 avss.n710 avss.n709 141.554
R1720 avss.n700 avss.n149 141.554
R1721 avss.n156 avss.n150 141.554
R1722 avss.n152 avss.n150 141.554
R1723 avss.n701 avss.n700 141.554
R1724 avss.n681 avss.n673 141.554
R1725 avss.n686 avss.n685 141.554
R1726 avss.n685 avss.n672 141.554
R1727 avss.n681 avss.n680 141.554
R1728 avss.n666 avss.n663 141.554
R1729 avss.n661 avss.n131 141.554
R1730 avss.n715 avss.n131 141.554
R1731 avss.n667 avss.n666 141.554
R1732 avss.t44 avss.n289 119.891
R1733 avss.n602 avss.t73 119.891
R1734 avss.n301 avss.n272 118.047
R1735 avss.n580 avss.n579 117.334
R1736 avss.n576 avss.n575 117.334
R1737 avss.n392 avss.n391 117.334
R1738 avss.n402 avss.n401 117.334
R1739 avss.n415 avss.n383 117.334
R1740 avss.n412 avss.n411 117.334
R1741 avss.n609 avss.n257 117.334
R1742 avss.n454 avss.n453 117.334
R1743 avss.n567 avss.n566 117.334
R1744 avss.n563 avss.n562 117.334
R1745 avss.n426 avss.n368 117.334
R1746 avss.n423 avss.n422 117.334
R1747 avss.n620 avss.n243 117.334
R1748 avss.n617 avss.n616 117.334
R1749 avss.n306 avss.n305 117.334
R1750 avss.n481 avss.n479 117.334
R1751 avss.n652 avss.n651 117.334
R1752 avss.n494 avss.n493 117.334
R1753 avss.n507 avss.n506 117.334
R1754 avss.n553 avss.n552 117.334
R1755 avss.n549 avss.n548 117.334
R1756 avss.n518 avss.n517 117.334
R1757 avss.n628 avss.n627 117.334
R1758 avss.n631 avss.n229 117.334
R1759 avss.n285 avss.n284 117.334
R1760 avss.n221 avss.n220 117.334
R1761 avss.n210 avss.n209 117.334
R1762 avss.n198 avss.n197 117.334
R1763 avss.n640 avss.n187 117.334
R1764 avss.t147 avss.n317 110.832
R1765 avss.n537 avss.t131 103.657
R1766 avss.n182 avss.t190 103.657
R1767 avss.n310 avss.n249 101.447
R1768 avss.n599 avss.n314 100.894
R1769 avss.n312 avss.n266 100.894
R1770 avss.n340 avss.n339 100.894
R1771 avss.n346 avss.n345 100.894
R1772 avss.n291 avss.n276 100.894
R1773 avss.n296 avss.n278 100.894
R1774 avss.n461 avss.n460 100.894
R1775 avss.n463 avss.n445 100.894
R1776 avss.n532 avss.n527 100.894
R1777 avss.n535 avss.n534 100.894
R1778 avss.n645 avss.n175 100.894
R1779 avss.n179 avss.n178 100.894
R1780 avss.n640 avss.n639 97.5005
R1781 avss.n639 avss.n167 97.5005
R1782 avss.n190 avss.n189 97.5005
R1783 avss.n637 avss.n190 97.5005
R1784 avss.n220 avss.n219 97.5005
R1785 avss.n219 avss.n161 97.5005
R1786 avss.n223 avss.n222 97.5005
R1787 avss.n224 avss.n223 97.5005
R1788 avss.n653 avss.n652 97.5005
R1789 avss.n654 avss.n653 97.5005
R1790 avss.n650 avss.n649 97.5005
R1791 avss.n649 avss.n648 97.5005
R1792 avss.n209 avss.n207 97.5005
R1793 avss.n207 avss.n206 97.5005
R1794 avss.n212 avss.n211 97.5005
R1795 avss.n213 avss.n212 97.5005
R1796 avss.n507 avss.n497 97.5005
R1797 avss.n502 avss.n497 97.5005
R1798 avss.n499 avss.n498 97.5005
R1799 avss.n503 avss.n499 97.5005
R1800 avss.n566 avss.n360 97.5005
R1801 avss.n430 avss.n360 97.5005
R1802 avss.n569 avss.n568 97.5005
R1803 avss.n570 avss.n569 97.5005
R1804 avss.n576 avss.n353 97.5005
R1805 avss.n572 avss.n353 97.5005
R1806 avss.n355 avss.n354 97.5005
R1807 avss.n355 avss.n318 97.5005
R1808 avss.n482 avss.n481 97.5005
R1809 avss.n483 avss.n482 97.5005
R1810 avss.n478 avss.n477 97.5005
R1811 avss.n477 avss.n476 97.5005
R1812 avss.n197 avss.n196 97.5005
R1813 avss.n196 avss.n195 97.5005
R1814 avss.n200 avss.n199 97.5005
R1815 avss.n201 avss.n200 97.5005
R1816 avss.n549 avss.n522 97.5005
R1817 avss.n544 avss.n522 97.5005
R1818 avss.n524 avss.n523 97.5005
R1819 avss.n545 avss.n524 97.5005
R1820 avss.n427 avss.n426 97.5005
R1821 avss.n428 avss.n427 97.5005
R1822 avss.n375 avss.n374 97.5005
R1823 avss.n376 avss.n375 97.5005
R1824 avss.n402 avss.n395 97.5005
R1825 avss.n398 avss.n395 97.5005
R1826 avss.n397 avss.n396 97.5005
R1827 avss.n397 avss.n319 97.5005
R1828 avss.n628 avss.n231 97.5005
R1829 avss.n234 avss.n231 97.5005
R1830 avss.n233 avss.n232 97.5005
R1831 avss.n624 avss.n233 97.5005
R1832 avss.n621 avss.n620 97.5005
R1833 avss.n622 avss.n621 97.5005
R1834 avss.n251 avss.n250 97.5005
R1835 avss.n252 avss.n251 97.5005
R1836 avss.n412 avss.n405 97.5005
R1837 avss.n408 avss.n405 97.5005
R1838 avss.n407 avss.n406 97.5005
R1839 avss.n407 avss.n320 97.5005
R1840 avss.n284 avss.n283 97.5005
R1841 avss.n283 avss.n225 97.5005
R1842 avss.n287 avss.n286 97.5005
R1843 avss.n288 avss.n287 97.5005
R1844 avss.n305 avss.n303 97.5005
R1845 avss.n303 avss.n302 97.5005
R1846 avss.n308 avss.n307 97.5005
R1847 avss.n309 avss.n308 97.5005
R1848 avss.n606 avss.n259 97.5005
R1849 avss.n264 avss.n259 97.5005
R1850 avss.n316 avss.n315 97.5005
R1851 avss.n593 avss.n316 97.5005
R1852 avss.n632 avss.n631 97.5005
R1853 avss.n633 avss.n632 97.5005
R1854 avss.n237 avss.n236 97.5005
R1855 avss.n238 avss.n237 97.5005
R1856 avss.n617 avss.n245 97.5005
R1857 avss.n248 avss.n245 97.5005
R1858 avss.n247 avss.n246 97.5005
R1859 avss.n613 avss.n247 97.5005
R1860 avss.n610 avss.n609 97.5005
R1861 avss.n611 avss.n610 97.5005
R1862 avss.n322 avss.n321 97.5005
R1863 avss.n323 avss.n322 97.5005
R1864 avss.n518 avss.n510 97.5005
R1865 avss.n513 avss.n510 97.5005
R1866 avss.n512 avss.n511 97.5005
R1867 avss.n514 avss.n512 97.5005
R1868 avss.n423 avss.n370 97.5005
R1869 avss.n373 avss.n370 97.5005
R1870 avss.n372 avss.n371 97.5005
R1871 avss.n419 avss.n372 97.5005
R1872 avss.n416 avss.n415 97.5005
R1873 avss.n417 avss.n416 97.5005
R1874 avss.n382 avss.n381 97.5005
R1875 avss.n381 avss.n324 97.5005
R1876 avss.n552 avss.n435 97.5005
R1877 avss.n500 avss.n435 97.5005
R1878 avss.n555 avss.n554 97.5005
R1879 avss.n556 avss.n555 97.5005
R1880 avss.n563 avss.n362 97.5005
R1881 avss.n558 avss.n362 97.5005
R1882 avss.n364 avss.n363 97.5005
R1883 avss.n559 avss.n364 97.5005
R1884 avss.n392 avss.n385 97.5005
R1885 avss.n388 avss.n385 97.5005
R1886 avss.n387 avss.n386 97.5005
R1887 avss.n387 avss.n325 97.5005
R1888 avss.n494 avss.n437 97.5005
R1889 avss.n440 avss.n437 97.5005
R1890 avss.n439 avss.n438 97.5005
R1891 avss.n490 avss.n439 97.5005
R1892 avss.n454 avss.n447 97.5005
R1893 avss.n447 avss.n441 97.5005
R1894 avss.n449 avss.n448 97.5005
R1895 avss.n450 avss.n449 97.5005
R1896 avss.n579 avss.n330 97.5005
R1897 avss.n330 avss.n329 97.5005
R1898 avss.n582 avss.n581 97.5005
R1899 avss.n583 avss.n582 97.5005
R1900 avss.t80 avss.n119 97.3856
R1901 avss.t80 avss.n121 97.3856
R1902 avss.n594 avss.n261 95.7798
R1903 avss.n634 avss.n225 87.6132
R1904 avss.n593 avss.n592 87.6132
R1905 avss.n636 avss.t131 83.1239
R1906 avss.n636 avss.t141 80.8829
R1907 avss.n541 avss.n527 72.1417
R1908 avss.n539 avss.n535 72.1417
R1909 avss.n645 avss.n644 68.4924
R1910 avss.n184 avss.n179 68.4924
R1911 avss.n339 avss.n332 67.468
R1912 avss.n346 avss.n331 67.468
R1913 avss.n299 avss.n276 67.468
R1914 avss.n297 avss.n296 67.468
R1915 avss.n460 avss.n457 67.468
R1916 avss.n470 avss.n445 67.468
R1917 avss.n668 avss.n667 65.0005
R1918 avss.n694 avss.n668 65.0005
R1919 avss.n661 avss.n138 65.0005
R1920 avss.n713 avss.n138 65.0005
R1921 avss.n663 avss.n160 65.0005
R1922 avss.n694 avss.n160 65.0005
R1923 avss.n715 avss.n714 65.0005
R1924 avss.n714 avss.n713 65.0005
R1925 avss.n687 avss.n686 65.0005
R1926 avss.n694 avss.n687 65.0005
R1927 avss.n673 avss.n139 65.0005
R1928 avss.n713 avss.n139 65.0005
R1929 avss.n672 avss.n159 65.0005
R1930 avss.n694 avss.n159 65.0005
R1931 avss.n680 avss.n136 65.0005
R1932 avss.n713 avss.n136 65.0005
R1933 avss.n695 avss.n156 65.0005
R1934 avss.n695 avss.n694 65.0005
R1935 avss.n149 avss.n140 65.0005
R1936 avss.n713 avss.n140 65.0005
R1937 avss.n153 avss.n152 65.0005
R1938 avss.n694 avss.n153 65.0005
R1939 avss.n701 avss.n135 65.0005
R1940 avss.n713 avss.n135 65.0005
R1941 avss.n693 avss.n692 65.0005
R1942 avss.n694 avss.n693 65.0005
R1943 avss.n712 avss.n711 65.0005
R1944 avss.n713 avss.n712 65.0005
R1945 avss.n690 avss.n158 65.0005
R1946 avss.n694 avss.n158 65.0005
R1947 avss.n709 avss.n134 65.0005
R1948 avss.n713 avss.n134 65.0005
R1949 avss.n737 avss.n111 62.759
R1950 avss.n730 avss.n116 61.5669
R1951 avss.n713 avss.n137 59.8963
R1952 avss.n731 avss.n730 59.0984
R1953 avss.n647 avss.t190 55.4161
R1954 avss.n647 avss.t161 53.9221
R1955 avss.n662 avss.n659 53.1823
R1956 avss.n659 avss.t31 53.1823
R1957 avss.n665 avss.n664 53.1823
R1958 avss.n664 avss.t31 53.1823
R1959 avss.n671 avss.n669 53.1823
R1960 avss.n669 avss.t31 53.1823
R1961 avss.n684 avss.n683 53.1823
R1962 avss.n683 avss.t31 53.1823
R1963 avss.n675 avss.n674 53.1823
R1964 avss.n674 avss.t31 53.1823
R1965 avss.n155 avss.n154 53.1823
R1966 avss.n154 avss.t31 53.1823
R1967 avss.n699 avss.n698 53.1823
R1968 avss.n698 avss.t31 53.1823
R1969 avss.n151 avss.n148 53.1823
R1970 avss.n151 avss.t31 53.1823
R1971 avss.n143 avss.n141 53.1823
R1972 avss.n141 avss.t31 53.1823
R1973 avss.n688 avss.n144 53.1823
R1974 avss.n688 avss.t31 53.1823
R1975 avss.n157 avss.n145 53.1823
R1976 avss.n157 avss.t31 53.1823
R1977 avss.n133 avss.n130 53.1823
R1978 avss.n657 avss.n133 53.1823
R1979 avss.n188 avss.n186 53.1823
R1980 avss.t25 avss.n188 53.1823
R1981 avss.n638 avss.n187 53.1823
R1982 avss.n638 avss.t25 53.1823
R1983 avss.n218 avss.n216 53.1823
R1984 avss.n216 avss.t60 53.1823
R1985 avss.n221 avss.n217 53.1823
R1986 avss.n217 avss.t60 53.1823
R1987 avss.n165 avss.n163 53.1823
R1988 avss.n163 avss.t41 53.1823
R1989 avss.n651 avss.n164 53.1823
R1990 avss.n164 avss.t41 53.1823
R1991 avss.n205 avss.n203 53.1823
R1992 avss.n203 avss.t26 53.1823
R1993 avss.n210 avss.n204 53.1823
R1994 avss.n204 avss.t26 53.1823
R1995 avss.n504 avss.n496 53.1823
R1996 avss.t217 avss.n504 53.1823
R1997 avss.n506 avss.n505 53.1823
R1998 avss.n505 avss.t217 53.1823
R1999 avss.n359 avss.n357 53.1823
R2000 avss.n357 avss.t148 53.1823
R2001 avss.n567 avss.n358 53.1823
R2002 avss.n358 avss.t148 53.1823
R2003 avss.n573 avss.n352 53.1823
R2004 avss.t157 avss.n573 53.1823
R2005 avss.n575 avss.n574 53.1823
R2006 avss.n574 avss.t157 53.1823
R2007 avss.n475 avss.n473 53.1823
R2008 avss.n473 avss.t246 53.1823
R2009 avss.n479 avss.n474 53.1823
R2010 avss.n474 avss.t246 53.1823
R2011 avss.n194 avss.n192 53.1823
R2012 avss.n192 avss.t254 53.1823
R2013 avss.n198 avss.n193 53.1823
R2014 avss.n193 avss.t254 53.1823
R2015 avss.n546 avss.n521 53.1823
R2016 avss.t216 avss.n546 53.1823
R2017 avss.n548 avss.n547 53.1823
R2018 avss.n547 avss.t216 53.1823
R2019 avss.n367 avss.n365 53.1823
R2020 avss.n365 avss.t136 53.1823
R2021 avss.n368 avss.n366 53.1823
R2022 avss.n366 avss.t136 53.1823
R2023 avss.n399 avss.n394 53.1823
R2024 avss.t191 avss.n399 53.1823
R2025 avss.n401 avss.n400 53.1823
R2026 avss.n400 avss.t191 53.1823
R2027 avss.n625 avss.n230 53.1823
R2028 avss.t214 avss.n625 53.1823
R2029 avss.n627 avss.n626 53.1823
R2030 avss.n626 avss.t214 53.1823
R2031 avss.n242 avss.n240 53.1823
R2032 avss.n240 avss.t101 53.1823
R2033 avss.n243 avss.n241 53.1823
R2034 avss.n241 avss.t101 53.1823
R2035 avss.n409 avss.n404 53.1823
R2036 avss.t30 avss.n409 53.1823
R2037 avss.n411 avss.n410 53.1823
R2038 avss.n410 avss.t30 53.1823
R2039 avss.n282 avss.n280 53.1823
R2040 avss.n280 avss.t215 53.1823
R2041 avss.n285 avss.n281 53.1823
R2042 avss.n281 avss.t215 53.1823
R2043 avss.n271 avss.n269 53.1823
R2044 avss.n269 avss.t158 53.1823
R2045 avss.n306 avss.n270 53.1823
R2046 avss.n270 avss.t158 53.1823
R2047 avss.n597 avss.n596 53.1823
R2048 avss.n596 avss.t61 53.1823
R2049 avss.n595 avss.n594 53.1823
R2050 avss.t61 avss.n595 53.1823
R2051 avss.n228 avss.n226 53.1823
R2052 avss.n226 avss.t187 53.1823
R2053 avss.n229 avss.n227 53.1823
R2054 avss.n227 avss.t187 53.1823
R2055 avss.n614 avss.n244 53.1823
R2056 avss.t197 avss.n614 53.1823
R2057 avss.n616 avss.n615 53.1823
R2058 avss.n615 avss.t197 53.1823
R2059 avss.n256 avss.n254 53.1823
R2060 avss.n254 avss.t151 53.1823
R2061 avss.n257 avss.n255 53.1823
R2062 avss.n255 avss.t151 53.1823
R2063 avss.n515 avss.n509 53.1823
R2064 avss.t112 avss.n515 53.1823
R2065 avss.n517 avss.n516 53.1823
R2066 avss.n516 avss.t112 53.1823
R2067 avss.n420 avss.n369 53.1823
R2068 avss.t239 avss.n420 53.1823
R2069 avss.n422 avss.n421 53.1823
R2070 avss.n421 avss.t239 53.1823
R2071 avss.n380 avss.n378 53.1823
R2072 avss.n378 avss.t47 53.1823
R2073 avss.n383 avss.n379 53.1823
R2074 avss.n379 avss.t47 53.1823
R2075 avss.n434 avss.n432 53.1823
R2076 avss.n432 avss.t188 53.1823
R2077 avss.n553 avss.n433 53.1823
R2078 avss.n433 avss.t188 53.1823
R2079 avss.n560 avss.n361 53.1823
R2080 avss.t182 avss.n560 53.1823
R2081 avss.n562 avss.n561 53.1823
R2082 avss.n561 avss.t182 53.1823
R2083 avss.n389 avss.n384 53.1823
R2084 avss.t29 avss.n389 53.1823
R2085 avss.n391 avss.n390 53.1823
R2086 avss.n390 avss.t29 53.1823
R2087 avss.n491 avss.n436 53.1823
R2088 avss.t186 avss.n491 53.1823
R2089 avss.n493 avss.n492 53.1823
R2090 avss.n492 avss.t186 53.1823
R2091 avss.n451 avss.n446 53.1823
R2092 avss.t57 avss.n451 53.1823
R2093 avss.n453 avss.n452 53.1823
R2094 avss.n452 avss.t57 53.1823
R2095 avss.n328 avss.n326 53.1823
R2096 avss.n326 avss.t196 53.1823
R2097 avss.n580 avss.n327 53.1823
R2098 avss.n327 avss.t196 53.1823
R2099 avss.n730 avss.n729 53.1823
R2100 avss.n729 avss.t80 53.1823
R2101 avss.n728 avss.n727 53.1823
R2102 avss.t80 avss.n728 53.1823
R2103 avss.n314 avss.n313 51.9534
R2104 avss.n313 avss.n312 51.9534
R2105 avss.n345 avss.n333 51.9534
R2106 avss.n340 avss.n333 51.9534
R2107 avss.n291 avss.n290 51.9534
R2108 avss.n290 avss.n278 51.9534
R2109 avss.n463 avss.n458 51.9534
R2110 avss.n461 avss.n458 51.9534
R2111 avss.n533 avss.n532 51.9534
R2112 avss.n534 avss.n533 51.9534
R2113 avss.n177 avss.n175 51.9534
R2114 avss.n178 avss.n177 51.9534
R2115 avss.n599 avss.n598 50.6259
R2116 avss.n313 avss.n260 48.9417
R2117 avss.n349 avss.n333 48.9417
R2118 avss.n290 avss.n277 48.9417
R2119 avss.n468 avss.n458 48.9417
R2120 avss.n533 avss.n528 48.9417
R2121 avss.n177 avss.n176 48.9417
R2122 avss.n118 avss.n115 48.7505
R2123 avss.n121 avss.n118 48.7505
R2124 avss.n123 avss.n117 48.7505
R2125 avss.n119 avss.n117 48.7505
R2126 avss.n266 avss.n261 43.6169
R2127 avss.n605 avss.n260 42.5417
R2128 avss.n350 avss.n349 42.5417
R2129 avss.n298 avss.n277 42.5417
R2130 avss.n469 avss.n468 42.5417
R2131 avss.n540 avss.n528 42.5417
R2132 avss.n643 avss.n176 42.5417
R2133 avss.n146 avss.t90 41.586
R2134 avss.n147 avss.t142 41.586
R2135 avss.n676 avss.t66 41.586
R2136 avss.n129 avss.t238 41.586
R2137 avss.n146 avss.t185 40.9588
R2138 avss.n147 avss.t32 40.9588
R2139 avss.n676 avss.t54 40.9588
R2140 avss.n129 avss.t247 40.9588
R2141 avss.n731 avss.n115 32.2212
R2142 avss.n589 avss.n122 31.0458
R2143 avss.n541 avss.n540 31.0005
R2144 avss.n540 avss.n539 31.0005
R2145 avss.n725 avss.t81 30.1756
R2146 avss.n589 avss.n588 29.7453
R2147 avss.n591 avss.t152 27.3441
R2148 avss.n585 avss.t152 27.3441
R2149 avss.n644 avss.n643 27.1786
R2150 avss.n643 avss.n184 27.1786
R2151 avss.n115 avss.n111 27.1769
R2152 avss.n350 avss.n331 26.1058
R2153 avss.n350 avss.n332 26.1058
R2154 avss.n299 avss.n298 26.1058
R2155 avss.n298 avss.n297 26.1058
R2156 avss.n470 avss.n469 26.1058
R2157 avss.n469 avss.n457 26.1058
R2158 avss.n585 avss.n119 24.3994
R2159 avss.n121 avss.n120 23.558
R2160 avss.n658 avss.t31 19.4289
R2161 avss.t73 avss.n249 18.4453
R2162 avss.n726 avss.n123 16.7152
R2163 avss.n737 avss.n736 11.7731
R2164 avss.n489 avss.t189 11.0836
R2165 avss.n123 avss.n116 10.9042
R2166 avss.n105 avss.t83 10.7251
R2167 avss.n4 avss.t220 10.6793
R2168 avss.n107 avss.t9 10.5739
R2169 avss.n109 avss.t105 10.5739
R2170 avss.n1 avss.t28 10.5739
R2171 avss.n3 avss.t221 10.5739
R2172 avss.n58 avss.t223 10.5739
R2173 avss.n57 avss.t181 10.5739
R2174 avss.n55 avss.t167 10.5739
R2175 avss.n53 avss.t34 10.5739
R2176 avss.n51 avss.t165 10.5739
R2177 avss.n50 avss.t144 10.5739
R2178 avss.n49 avss.t72 10.5739
R2179 avss.n48 avss.t156 10.5739
R2180 avss.n47 avss.t116 10.5739
R2181 avss.n46 avss.t79 10.5739
R2182 avss.n45 avss.t150 10.5739
R2183 avss.n44 avss.t107 10.5739
R2184 avss.n43 avss.t207 10.5739
R2185 avss.n42 avss.t43 10.5739
R2186 avss.n41 avss.t111 10.5739
R2187 avss.n40 avss.t175 10.5739
R2188 avss.n39 avss.t124 10.5739
R2189 avss.n38 avss.t211 10.5739
R2190 avss.n37 avss.t193 10.5739
R2191 avss.n36 avss.t16 10.5739
R2192 avss.n35 avss.t118 10.5739
R2193 avss.n34 avss.t233 10.5739
R2194 avss.n33 avss.t179 10.5739
R2195 avss.n32 avss.t65 10.5739
R2196 avss.n31 avss.t209 10.5739
R2197 avss.n30 avss.t225 10.5739
R2198 avss.n29 avss.t103 10.5739
R2199 avss.n28 avss.t96 10.5739
R2200 avss.n27 avss.t199 10.5739
R2201 avss.n26 avss.t177 10.5739
R2202 avss.n25 avss.t38 10.5739
R2203 avss.n24 avss.t201 10.5739
R2204 avss.n23 avss.t243 10.5739
R2205 avss.n22 avss.t130 10.5739
R2206 avss.n21 avss.t75 10.5739
R2207 avss.n20 avss.t195 10.5739
R2208 avss.n19 avss.t227 10.5739
R2209 avss.n18 avss.t63 10.5739
R2210 avss.n17 avss.t53 10.5739
R2211 avss.n16 avss.t51 10.5739
R2212 avss.n15 avss.t77 10.5739
R2213 avss.n14 avss.t122 10.5739
R2214 avss.n13 avss.t46 10.5739
R2215 avss.n12 avss.t163 10.5739
R2216 avss.n11 avss.t138 10.5739
R2217 avss.n10 avss.t70 10.5739
R2218 avss.n9 avss.t92 10.5739
R2219 avss.n8 avss.t128 10.5739
R2220 avss.n7 avss.t109 10.5739
R2221 avss.n6 avss.t24 10.5739
R2222 avss.n5 avss.t20 10.5739
R2223 avss.n59 avss.t68 10.5739
R2224 avss.n60 avss.t235 10.5739
R2225 avss.n61 avss.t253 10.5739
R2226 avss.n62 avss.t36 10.5739
R2227 avss.n63 avss.t94 10.5739
R2228 avss.n64 avss.t154 10.5739
R2229 avss.n65 avss.t171 10.5739
R2230 avss.n66 avss.t126 10.5739
R2231 avss.n67 avss.t56 10.5739
R2232 avss.n68 avss.t98 10.5739
R2233 avss.n69 avss.t256 10.5739
R2234 avss.n70 avss.t140 10.5739
R2235 avss.n71 avss.t49 10.5739
R2236 avss.n72 avss.t133 10.5739
R2237 avss.n73 avss.t231 10.5739
R2238 avss.n74 avss.t173 10.5739
R2239 avss.n75 avss.t169 10.5739
R2240 avss.n76 avss.t59 10.5739
R2241 avss.n77 avss.t114 10.5739
R2242 avss.n78 avss.t87 10.5739
R2243 avss.n79 avss.t7 10.5739
R2244 avss.n80 avss.t241 10.5739
R2245 avss.n81 avss.t205 10.5739
R2246 avss.n82 avss.t85 10.5739
R2247 avss.n83 avss.t251 10.5739
R2248 avss.n84 avss.t2 10.5739
R2249 avss.n85 avss.t219 10.5739
R2250 avss.n86 avss.t184 10.5739
R2251 avss.n87 avss.t237 10.5739
R2252 avss.n88 avss.t146 10.5739
R2253 avss.n89 avss.t203 10.5739
R2254 avss.n90 avss.t245 10.5739
R2255 avss.n91 avss.t22 10.5739
R2256 avss.n92 avss.t89 10.5739
R2257 avss.n93 avss.t12 10.5739
R2258 avss.n94 avss.t4 10.5739
R2259 avss.n95 avss.t40 10.5739
R2260 avss.n96 avss.t120 10.5739
R2261 avss.n97 avss.t258 10.5739
R2262 avss.n98 avss.t135 10.5739
R2263 avss.n99 avss.t18 10.5739
R2264 avss.n100 avss.t100 10.5739
R2265 avss.n101 avss.t229 10.5739
R2266 avss.n102 avss.t213 10.5739
R2267 avss.n103 avss.t160 10.5739
R2268 avss.n104 avss.t249 10.5739
R2269 avss.n5 avss.t19 10.5285
R2270 avss.n6 avss.t23 10.5285
R2271 avss.n7 avss.t108 10.5285
R2272 avss.n8 avss.t127 10.5285
R2273 avss.n9 avss.t91 10.5285
R2274 avss.n10 avss.t69 10.5285
R2275 avss.n11 avss.t137 10.5285
R2276 avss.n12 avss.t162 10.5285
R2277 avss.n13 avss.t45 10.5285
R2278 avss.n14 avss.t121 10.5285
R2279 avss.n15 avss.t76 10.5285
R2280 avss.n16 avss.t50 10.5285
R2281 avss.n17 avss.t52 10.5285
R2282 avss.n18 avss.t62 10.5285
R2283 avss.n19 avss.t226 10.5285
R2284 avss.n20 avss.t194 10.5285
R2285 avss.n21 avss.t74 10.5285
R2286 avss.n22 avss.t129 10.5285
R2287 avss.n23 avss.t242 10.5285
R2288 avss.n24 avss.t200 10.5285
R2289 avss.n25 avss.t37 10.5285
R2290 avss.n26 avss.t176 10.5285
R2291 avss.n27 avss.t198 10.5285
R2292 avss.n28 avss.t95 10.5285
R2293 avss.n29 avss.t102 10.5285
R2294 avss.n30 avss.t224 10.5285
R2295 avss.n31 avss.t208 10.5285
R2296 avss.n32 avss.t64 10.5285
R2297 avss.n33 avss.t178 10.5285
R2298 avss.n34 avss.t232 10.5285
R2299 avss.n35 avss.t117 10.5285
R2300 avss.n36 avss.t15 10.5285
R2301 avss.n37 avss.t192 10.5285
R2302 avss.n38 avss.t210 10.5285
R2303 avss.n39 avss.t123 10.5285
R2304 avss.n40 avss.t174 10.5285
R2305 avss.n41 avss.t110 10.5285
R2306 avss.n42 avss.t42 10.5285
R2307 avss.n43 avss.t206 10.5285
R2308 avss.n44 avss.t106 10.5285
R2309 avss.n45 avss.t149 10.5285
R2310 avss.n46 avss.t78 10.5285
R2311 avss.n47 avss.t115 10.5285
R2312 avss.n48 avss.t155 10.5285
R2313 avss.n49 avss.t71 10.5285
R2314 avss.n50 avss.t143 10.5285
R2315 avss.n51 avss.t164 10.5285
R2316 avss.n52 avss.t33 10.5285
R2317 avss.n54 avss.t166 10.5285
R2318 avss.n56 avss.t180 10.5285
R2319 avss.n104 avss.t248 10.5285
R2320 avss.n103 avss.t159 10.5285
R2321 avss.n102 avss.t212 10.5285
R2322 avss.n101 avss.t228 10.5285
R2323 avss.n100 avss.t99 10.5285
R2324 avss.n99 avss.t17 10.5285
R2325 avss.n98 avss.t134 10.5285
R2326 avss.n97 avss.t257 10.5285
R2327 avss.n96 avss.t119 10.5285
R2328 avss.n95 avss.t39 10.5285
R2329 avss.n94 avss.t3 10.5285
R2330 avss.n93 avss.t11 10.5285
R2331 avss.n92 avss.t88 10.5285
R2332 avss.n91 avss.t21 10.5285
R2333 avss.n90 avss.t244 10.5285
R2334 avss.n89 avss.t202 10.5285
R2335 avss.n88 avss.t145 10.5285
R2336 avss.n87 avss.t236 10.5285
R2337 avss.n86 avss.t183 10.5285
R2338 avss.n85 avss.t218 10.5285
R2339 avss.n84 avss.t1 10.5285
R2340 avss.n83 avss.t250 10.5285
R2341 avss.n82 avss.t84 10.5285
R2342 avss.n81 avss.t204 10.5285
R2343 avss.n80 avss.t240 10.5285
R2344 avss.n79 avss.t6 10.5285
R2345 avss.n78 avss.t86 10.5285
R2346 avss.n77 avss.t113 10.5285
R2347 avss.n76 avss.t58 10.5285
R2348 avss.n75 avss.t168 10.5285
R2349 avss.n74 avss.t172 10.5285
R2350 avss.n73 avss.t230 10.5285
R2351 avss.n72 avss.t132 10.5285
R2352 avss.n71 avss.t48 10.5285
R2353 avss.n70 avss.t139 10.5285
R2354 avss.n69 avss.t255 10.5285
R2355 avss.n68 avss.t97 10.5285
R2356 avss.n67 avss.t55 10.5285
R2357 avss.n66 avss.t125 10.5285
R2358 avss.n65 avss.t170 10.5285
R2359 avss.n64 avss.t153 10.5285
R2360 avss.n63 avss.t93 10.5285
R2361 avss.n62 avss.t35 10.5285
R2362 avss.n61 avss.t252 10.5285
R2363 avss.n60 avss.t234 10.5285
R2364 avss.n59 avss.t67 10.5285
R2365 avss.n58 avss.t222 10.5285
R2366 avss.n2 avss.t27 10.5285
R2367 avss.n0 avss.t104 10.5285
R2368 avss.n108 avss.t8 10.5285
R2369 avss.n106 avss.t82 10.5285
R2370 avss.n592 avss.n591 10.3069
R2371 avss.n605 avss.n604 7.9365
R2372 avss.n727 avss.n726 7.29749
R2373 avss.n606 avss.n258 7.2709
R2374 avss.n604 avss.n261 6.4005
R2375 avss.n588 avss.n116 5.91288
R2376 avss.n727 avss.n111 5.86875
R2377 avss.n720 avss.n127 5.34317
R2378 avss.n598 avss.n258 5.1205
R2379 avss.n721 avss.n126 3.60826
R2380 avss.n723 avss.n124 3.46074
R2381 avss.n722 avss.n125 3.42275
R2382 avss.n736 avss.n735 2.91095
R2383 avss.n735 avss.t10 2.91095
R2384 avss.n734 avss.n733 2.91095
R2385 avss.t10 avss.n734 2.91095
R2386 avss.n652 avss 2.78541
R2387 avss.n208 avss 2.23541
R2388 avss.n641 avss 2.23541
R2389 avss.n720 avss.n719 2.20222
R2390 avss.n732 avss.n113 2.19151
R2391 avss.n120 avss.n113 2.19151
R2392 avss.n114 avss.n112 2.19151
R2393 avss.t44 avss.n272 1.84498
R2394 avss.n726 avss.n122 1.80664
R2395 avss.n607 avss.n606 1.5505
R2396 avss.n609 avss.n608 1.5505
R2397 avss.n413 avss.n412 1.5505
R2398 avss.n415 avss.n414 1.5505
R2399 avss.n403 avss.n402 1.5505
R2400 avss.n393 avss.n392 1.5505
R2401 avss.n577 avss.n576 1.5505
R2402 avss.n579 avss.n578 1.5505
R2403 avss.n305 avss.n304 1.5505
R2404 avss.n618 avss.n617 1.5505
R2405 avss.n620 avss.n619 1.5505
R2406 avss.n424 avss.n423 1.5505
R2407 avss.n426 avss.n425 1.5505
R2408 avss.n564 avss.n563 1.5505
R2409 avss.n566 avss.n565 1.5505
R2410 avss.n455 avss.n454 1.5505
R2411 avss.n481 avss.n480 1.5505
R2412 avss.n550 avss.n549 1.5505
R2413 avss.n552 avss.n551 1.5505
R2414 avss.n508 avss.n507 1.5505
R2415 avss.n495 avss.n494 1.5505
R2416 avss.n284 avss.n126 1.5505
R2417 avss.n631 avss.n630 1.5505
R2418 avss.n629 avss.n628 1.5505
R2419 avss.n519 avss.n518 1.5505
R2420 avss.n197 avss.n185 1.5505
R2421 avss.n209 avss.n208 1.5505
R2422 avss.n220 avss.n127 1.5505
R2423 avss.n641 avss.n640 1.5505
R2424 avss.n53 avss.n52 1.42736
R2425 avss.n55 avss.n54 1.42736
R2426 avss.n57 avss.n56 1.42736
R2427 avss.n2 avss.n1 1.42736
R2428 avss.n108 avss.n107 1.42736
R2429 avss.n706 avss.n705 1.37676
R2430 avss.n110 avss 1.34985
R2431 avss.n705 avss.n128 1.25238
R2432 avss.n719 avss.n128 1.25238
R2433 avss avss.n577 1.23541
R2434 avss.n393 avss 1.23541
R2435 avss.n403 avss 1.23541
R2436 avss.n414 avss 1.23541
R2437 avss avss.n413 1.23541
R2438 avss.n608 avss 1.23541
R2439 avss.n565 avss 1.23541
R2440 avss avss.n564 1.23541
R2441 avss.n425 avss 1.23541
R2442 avss avss.n424 1.23541
R2443 avss.n619 avss 1.23541
R2444 avss avss.n618 1.23541
R2445 avss.n480 avss 1.23541
R2446 avss.n495 avss 1.23541
R2447 avss.n508 avss 1.23541
R2448 avss.n551 avss 1.23541
R2449 avss avss.n550 1.23541
R2450 avss.n629 avss 1.23541
R2451 avss.n630 avss 1.23541
R2452 avss avss.n126 1.23541
R2453 avss.n208 avss 1.23541
R2454 avss avss.n185 1.23541
R2455 avss avss.n127 1.23541
R2456 avss.n605 avss.n124 1.163
R2457 avss.n351 avss.n350 1.163
R2458 avss.n298 avss.n125 1.163
R2459 avss.n469 avss.n456 1.163
R2460 avss.n540 avss.n520 1.163
R2461 avss.n643 avss.n642 1.163
R2462 avss avss.n519 1.11353
R2463 avss avss.n641 1.11353
R2464 avss avss.n607 1.10745
R2465 avss.n304 avss 1.07104
R2466 avss.n726 avss.n725 0.816777
R2467 avss.n578 avss.n351 0.74738
R2468 avss.n739 avss.n109 0.714152
R2469 avss.n739 avss.n0 0.713709
R2470 avss.n456 avss.n455 0.709387
R2471 avss.n606 avss.n605 0.6661
R2472 avss.n578 avss 0.5005
R2473 avss.n577 avss 0.5005
R2474 avss avss.n393 0.5005
R2475 avss avss.n403 0.5005
R2476 avss.n414 avss 0.5005
R2477 avss.n413 avss 0.5005
R2478 avss.n608 avss 0.5005
R2479 avss.n455 avss 0.5005
R2480 avss.n565 avss 0.5005
R2481 avss.n564 avss 0.5005
R2482 avss.n425 avss 0.5005
R2483 avss.n424 avss 0.5005
R2484 avss.n619 avss 0.5005
R2485 avss.n618 avss 0.5005
R2486 avss.n480 avss 0.5005
R2487 avss avss.n495 0.5005
R2488 avss avss.n508 0.5005
R2489 avss.n551 avss 0.5005
R2490 avss.n519 avss 0.5005
R2491 avss avss.n629 0.5005
R2492 avss.n630 avss 0.5005
R2493 avss.n740 avss.n739 0.459809
R2494 avss.n708 avss.n707 0.388
R2495 avss.n703 avss.n702 0.388
R2496 avss.n679 avss.n678 0.388
R2497 avss.n717 avss.n716 0.388
R2498 avss.n738 avss.n110 0.377227
R2499 avss.n706 avss.n146 0.329037
R2500 avss.n704 avss.n147 0.329037
R2501 avss.n677 avss.n676 0.329037
R2502 avss.n718 avss.n129 0.329037
R2503 avss.n707 avss 0.301379
R2504 avss.n703 avss 0.301379
R2505 avss.n678 avss 0.301379
R2506 avss.n717 avss 0.301379
R2507 avss.n550 avss.n520 0.274922
R2508 avss.n642 avss.n185 0.274922
R2509 avss.n707 avss.n706 0.258038
R2510 avss.n704 avss.n703 0.258038
R2511 avss.n678 avss.n677 0.258038
R2512 avss.n718 avss.n717 0.258038
R2513 avss.n54 avss.n53 0.238532
R2514 avss.n56 avss.n55 0.238532
R2515 avss.n3 avss.n2 0.238532
R2516 avss.n1 avss.n0 0.238532
R2517 avss.n109 avss.n108 0.238532
R2518 avss.n107 avss.n106 0.238532
R2519 avss.n351 avss 0.221517
R2520 avss.n724 avss.n110 0.191699
R2521 avss.n456 avss 0.183525
R2522 avss.n722 avss.n721 0.161722
R2523 avss.n721 avss.n720 0.160761
R2524 avss.n723 avss.n722 0.157495
R2525 avss.n4 avss.n3 0.151652
R2526 avss.n106 avss.n105 0.151209
R2527 avss.n52 avss.n51 0.142787
R2528 avss.n58 avss.n57 0.142344
R2529 avss.n740 avss 0.136236
R2530 avss.n724 avss.n723 0.133859
R2531 avss.n705 avss.n704 0.124872
R2532 avss.n677 avss.n128 0.124872
R2533 avss.n719 avss.n718 0.124872
R2534 avss avss.n740 0.0871641
R2535 avss.n739 avss.n738 0.0830826
R2536 avss.n708 avss.n145 0.0554356
R2537 avss.n702 avss.n148 0.0554356
R2538 avss.n679 avss.n675 0.0554356
R2539 avss.n716 avss.n130 0.0554356
R2540 avss.n51 avss.n50 0.0429147
R2541 avss.n50 avss.n49 0.0429147
R2542 avss.n49 avss.n48 0.0429147
R2543 avss.n48 avss.n47 0.0429147
R2544 avss.n47 avss.n46 0.0429147
R2545 avss.n46 avss.n45 0.0429147
R2546 avss.n45 avss.n44 0.0429147
R2547 avss.n44 avss.n43 0.0429147
R2548 avss.n43 avss.n42 0.0429147
R2549 avss.n42 avss.n41 0.0429147
R2550 avss.n41 avss.n40 0.0429147
R2551 avss.n40 avss.n39 0.0429147
R2552 avss.n39 avss.n38 0.0429147
R2553 avss.n38 avss.n37 0.0429147
R2554 avss.n37 avss.n36 0.0429147
R2555 avss.n36 avss.n35 0.0429147
R2556 avss.n35 avss.n34 0.0429147
R2557 avss.n34 avss.n33 0.0429147
R2558 avss.n33 avss.n32 0.0429147
R2559 avss.n32 avss.n31 0.0429147
R2560 avss.n31 avss.n30 0.0429147
R2561 avss.n30 avss.n29 0.0429147
R2562 avss.n29 avss.n28 0.0429147
R2563 avss.n28 avss.n27 0.0429147
R2564 avss.n27 avss.n26 0.0429147
R2565 avss.n26 avss.n25 0.0429147
R2566 avss.n25 avss.n24 0.0429147
R2567 avss.n24 avss.n23 0.0429147
R2568 avss.n23 avss.n22 0.0429147
R2569 avss.n22 avss.n21 0.0429147
R2570 avss.n21 avss.n20 0.0429147
R2571 avss.n20 avss.n19 0.0429147
R2572 avss.n19 avss.n18 0.0429147
R2573 avss.n18 avss.n17 0.0429147
R2574 avss.n17 avss.n16 0.0429147
R2575 avss.n16 avss.n15 0.0429147
R2576 avss.n15 avss.n14 0.0429147
R2577 avss.n14 avss.n13 0.0429147
R2578 avss.n13 avss.n12 0.0429147
R2579 avss.n12 avss.n11 0.0429147
R2580 avss.n11 avss.n10 0.0429147
R2581 avss.n10 avss.n9 0.0429147
R2582 avss.n9 avss.n8 0.0429147
R2583 avss.n8 avss.n7 0.0429147
R2584 avss.n7 avss.n6 0.0429147
R2585 avss.n6 avss.n5 0.0429147
R2586 avss.n59 avss.n58 0.0429147
R2587 avss.n60 avss.n59 0.0429147
R2588 avss.n61 avss.n60 0.0429147
R2589 avss.n62 avss.n61 0.0429147
R2590 avss.n63 avss.n62 0.0429147
R2591 avss.n64 avss.n63 0.0429147
R2592 avss.n65 avss.n64 0.0429147
R2593 avss.n66 avss.n65 0.0429147
R2594 avss.n67 avss.n66 0.0429147
R2595 avss.n68 avss.n67 0.0429147
R2596 avss.n69 avss.n68 0.0429147
R2597 avss.n70 avss.n69 0.0429147
R2598 avss.n71 avss.n70 0.0429147
R2599 avss.n72 avss.n71 0.0429147
R2600 avss.n73 avss.n72 0.0429147
R2601 avss.n74 avss.n73 0.0429147
R2602 avss.n75 avss.n74 0.0429147
R2603 avss.n76 avss.n75 0.0429147
R2604 avss.n77 avss.n76 0.0429147
R2605 avss.n78 avss.n77 0.0429147
R2606 avss.n79 avss.n78 0.0429147
R2607 avss.n80 avss.n79 0.0429147
R2608 avss.n81 avss.n80 0.0429147
R2609 avss.n82 avss.n81 0.0429147
R2610 avss.n83 avss.n82 0.0429147
R2611 avss.n84 avss.n83 0.0429147
R2612 avss.n85 avss.n84 0.0429147
R2613 avss.n86 avss.n85 0.0429147
R2614 avss.n87 avss.n86 0.0429147
R2615 avss.n88 avss.n87 0.0429147
R2616 avss.n89 avss.n88 0.0429147
R2617 avss.n90 avss.n89 0.0429147
R2618 avss.n91 avss.n90 0.0429147
R2619 avss.n92 avss.n91 0.0429147
R2620 avss.n93 avss.n92 0.0429147
R2621 avss.n94 avss.n93 0.0429147
R2622 avss.n95 avss.n94 0.0429147
R2623 avss.n96 avss.n95 0.0429147
R2624 avss.n97 avss.n96 0.0429147
R2625 avss.n98 avss.n97 0.0429147
R2626 avss.n99 avss.n98 0.0429147
R2627 avss.n100 avss.n99 0.0429147
R2628 avss.n101 avss.n100 0.0429147
R2629 avss.n102 avss.n101 0.0429147
R2630 avss.n103 avss.n102 0.0429147
R2631 avss.n104 avss.n103 0.0429147
R2632 avss.n520 avss 0.0390514
R2633 avss.n642 avss 0.0390514
R2634 avss.n5 avss.n4 0.0270934
R2635 avss.n105 avss.n104 0.0270934
R2636 avss.n725 avss.n724 0.025588
R2637 avss.n607 avss.n124 0.00896354
R2638 avss.n738 avss.n737 0.00821144
R2639 avss.n304 avss.n125 0.00738559
R2640 multiplexer_0.vtrip_1_b.n0 multiplexer_0.vtrip_1_b.t0 41.0738
R2641 multiplexer_0.vtrip_1_b.n1 multiplexer_0.vtrip_1_b.n0 4.08093
R2642 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n13 0.521333
R2643 multiplexer_0.vtrip_1_b.n13 multiplexer_0.vtrip_1_b.n1 2.87169
R2644 multiplexer_0.vtrip_1_b.n13 multiplexer_0.vtrip_1_b.t6 33.8377
R2645 multiplexer_0.vtrip_1_b.t6 multiplexer_0.vtrip_1_b.n12 33.8377
R2646 multiplexer_0.vtrip_1_b.n12 multiplexer_0.vtrip_1_b.n11 17.2541
R2647 multiplexer_0.vtrip_1_b.n1 multiplexer_0.vtrip_1_b.n12 2.69901
R2648 multiplexer_0.vtrip_1_b.n9 multiplexer_0.vtrip_1_b.n10 0.315527
R2649 multiplexer_0.vtrip_1_b.n7 multiplexer_0.vtrip_1_b.n9 1.02307
R2650 multiplexer_0.vtrip_1_b.n5 multiplexer_0.vtrip_1_b.n7 1.02307
R2651 multiplexer_0.vtrip_1_b.n11 multiplexer_0.vtrip_1_b.n5 0.0551216
R2652 multiplexer_0.vtrip_1_b.n11 multiplexer_0.vtrip_1_b.n3 0.968446
R2653 multiplexer_0.vtrip_1_b.n10 multiplexer_0.vtrip_1_b.t2 99.1756
R2654 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n10 0.180561
R2655 multiplexer_0.vtrip_1_b.n3 multiplexer_0.vtrip_1_b.t4 99.4875
R2656 multiplexer_0.vtrip_1_b.n9 multiplexer_0.vtrip_1_b 2.77693
R2657 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n8 1.67907
R2658 multiplexer_0.vtrip_1_b.t8 multiplexer_0.vtrip_1_b.n8 16.8731
R2659 multiplexer_0.vtrip_1_b.n8 multiplexer_0.vtrip_1_b.t11 16.5088
R2660 multiplexer_0.vtrip_1_b.n7 multiplexer_0.vtrip_1_b 2.77693
R2661 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n6 1.67907
R2662 multiplexer_0.vtrip_1_b.t5 multiplexer_0.vtrip_1_b.n6 16.8731
R2663 multiplexer_0.vtrip_1_b.n6 multiplexer_0.vtrip_1_b.t7 16.5088
R2664 multiplexer_0.vtrip_1_b.n5 multiplexer_0.vtrip_1_b 2.77693
R2665 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n4 1.67907
R2666 multiplexer_0.vtrip_1_b.t12 multiplexer_0.vtrip_1_b.n4 16.8731
R2667 multiplexer_0.vtrip_1_b.n4 multiplexer_0.vtrip_1_b.t3 16.5088
R2668 multiplexer_0.vtrip_1_b.n3 multiplexer_0.vtrip_1_b 2.77693
R2669 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1_b.n2 1.67907
R2670 multiplexer_0.vtrip_1_b.t9 multiplexer_0.vtrip_1_b.n2 16.8731
R2671 multiplexer_0.vtrip_1_b.n2 multiplexer_0.vtrip_1_b.t10 16.5088
R2672 multiplexer_0.vtrip_1_b.n0 multiplexer_0.vtrip_1_b.t1 227.512
R2673 a_n15874_n447.t0 a_n15874_n447.t1 21.2567
R2674 a_n12654_n447.t0 a_n12654_n447.t1 21.34
R2675 a_n12118_12027.t0 a_n12118_12027.t1 21.2567
R2676 a_n8898_11649.t0 a_n8898_11649.t1 21.167
R2677 comp_hyst_0.net4.t0 comp_hyst_0.net4.n24 239.264
R2678 comp_hyst_0.net4.n23 comp_hyst_0.net4.n24 3.74168
R2679 comp_hyst_0.net4.n24 comp_hyst_0.net4.t12 9.62718
R2680 comp_hyst_0.net4.n3 comp_hyst_0.net4.n2 1.7055
R2681 comp_hyst_0.net4.n8 comp_hyst_0.net4.n7 1.7055
R2682 comp_hyst_0.net4.n23 comp_hyst_0.net4.n22 0.22541
R2683 comp_hyst_0.net4.n21 comp_hyst_0.net4.n23 0.20337
R2684 comp_hyst_0.net4.n13 comp_hyst_0.net4.n21 0.0768069
R2685 comp_hyst_0.net4.n12 comp_hyst_0.net4.n13 0.0948632
R2686 comp_hyst_0.net4.n3 comp_hyst_0.net4.n12 0.0950311
R2687 comp_hyst_0.net4.n8 comp_hyst_0.net4.n3 0.0472345
R2688 comp_hyst_0.net4.n1 comp_hyst_0.net4.n8 0.0950311
R2689 comp_hyst_0.net4.n0 comp_hyst_0.net4.n1 0.0908919
R2690 comp_hyst_0.net4 comp_hyst_0.net4.n0 0.0441783
R2691 comp_hyst_0.net4.n22 comp_hyst_0.net4.t8 85.3843
R2692 comp_hyst_0.net4.n22 comp_hyst_0.net4.t9 84.8697
R2693 comp_hyst_0.net4.n14 comp_hyst_0.net4.n16 12.7683
R2694 comp_hyst_0.net4.n21 comp_hyst_0.net4.n14 3.24613
R2695 comp_hyst_0.net4.n16 comp_hyst_0.net4.n15 0.3295
R2696 comp_hyst_0.net4.n17 comp_hyst_0.net4.n15 12.7689
R2697 comp_hyst_0.net4.n20 comp_hyst_0.net4.n17 1.66612
R2698 comp_hyst_0.net4.n2 comp_hyst_0.net4.n20 0.0663683
R2699 comp_hyst_0.net4.n7 comp_hyst_0.net4.n20 0.0663683
R2700 comp_hyst_0.net4.n14 comp_hyst_0.net4.n19 1.88237
R2701 comp_hyst_0.net4.n19 comp_hyst_0.net4.n18 0.3295
R2702 comp_hyst_0.net4.n17 comp_hyst_0.net4.n18 1.88299
R2703 comp_hyst_0.net4.n19 comp_hyst_0.net4.t7 231.423
R2704 comp_hyst_0.net4.n18 comp_hyst_0.net4.t5 231.423
R2705 comp_hyst_0.net4.n16 comp_hyst_0.net4.t6 231.423
R2706 comp_hyst_0.net4.n15 comp_hyst_0.net4.t10 231.423
R2707 comp_hyst_0.net4.n13 comp_hyst_0.net4.t11 8.12591
R2708 comp_hyst_0.net4.n12 comp_hyst_0.net4.n9 4.32456
R2709 comp_hyst_0.net4.n9 comp_hyst_0.net4.n10 2.00279
R2710 comp_hyst_0.net4.n11 comp_hyst_0.net4.n10 2.00279
R2711 comp_hyst_0.net4.n11 comp_hyst_0.net4.t1 11.9724
R2712 comp_hyst_0.net4.n9 comp_hyst_0.net4.t1 11.9724
R2713 comp_hyst_0.net4.n2 comp_hyst_0.net4.n11 2.4805
R2714 comp_hyst_0.net4.n10 comp_hyst_0.net4.t2 228.215
R2715 comp_hyst_0.net4.n7 comp_hyst_0.net4.n6 2.48206
R2716 comp_hyst_0.net4.n6 comp_hyst_0.net4.t3 11.9744
R2717 comp_hyst_0.net4.n6 comp_hyst_0.net4.n4 2.00084
R2718 comp_hyst_0.net4.n5 comp_hyst_0.net4.n4 2.00279
R2719 comp_hyst_0.net4.t3 comp_hyst_0.net4.n5 11.9724
R2720 comp_hyst_0.net4.n1 comp_hyst_0.net4.n5 4.32456
R2721 comp_hyst_0.net4.n4 comp_hyst_0.net4.t4 228.215
R2722 comp_hyst_0.net4.n0 comp_hyst_0.net4.t13 8.12988
R2723 dvdd.n534 dvdd.n98 6151.76
R2724 dvdd.n528 dvdd.n98 6151.76
R2725 dvdd.n528 dvdd.n57 6151.76
R2726 dvdd.n546 dvdd.n57 6151.76
R2727 dvdd.n546 dvdd.n71 6151.76
R2728 dvdd.n633 dvdd.n71 6151.76
R2729 dvdd.n533 dvdd.n99 6151.76
R2730 dvdd.n527 dvdd.n99 6151.76
R2731 dvdd.n527 dvdd.n58 6151.76
R2732 dvdd.n545 dvdd.n58 6151.76
R2733 dvdd.n545 dvdd.n72 6151.76
R2734 dvdd.n635 dvdd.n72 6151.76
R2735 dvdd.n622 dvdd.n94 6151.76
R2736 dvdd.n622 dvdd.n96 6151.76
R2737 dvdd.n96 dvdd.n59 6151.76
R2738 dvdd.n543 dvdd.n59 6151.76
R2739 dvdd.n543 dvdd.n73 6151.76
R2740 dvdd.n632 dvdd.n73 6151.76
R2741 dvdd.n621 dvdd.n101 6151.76
R2742 dvdd.n621 dvdd.n53 6151.76
R2743 dvdd.n659 dvdd.n53 6151.76
R2744 dvdd.n659 dvdd.n54 6151.76
R2745 dvdd.n653 dvdd.n54 6151.76
R2746 dvdd.n653 dvdd.n74 6151.76
R2747 dvdd.n111 dvdd.n100 6151.76
R2748 dvdd.n100 dvdd.n60 6151.76
R2749 dvdd.n658 dvdd.n60 6151.76
R2750 dvdd.n658 dvdd.n61 6151.76
R2751 dvdd.n654 dvdd.n61 6151.76
R2752 dvdd.n654 dvdd.n69 6151.76
R2753 dvdd.n589 dvdd.n268 4207.06
R2754 dvdd.n592 dvdd.n591 4207.06
R2755 dvdd.n227 dvdd.n139 3328.24
R2756 dvdd.n147 dvdd.n139 3328.24
R2757 dvdd.n242 dvdd.n132 3328.24
R2758 dvdd.n243 dvdd.n242 3328.24
R2759 dvdd.n169 dvdd.n138 3328.24
R2760 dvdd.n182 dvdd.n138 3328.24
R2761 dvdd.n201 dvdd.n137 3328.24
R2762 dvdd.n191 dvdd.n137 3328.24
R2763 dvdd.n170 dvdd.n136 3328.24
R2764 dvdd.n193 dvdd.n136 3328.24
R2765 dvdd.n241 dvdd.n141 3328.24
R2766 dvdd.n241 dvdd.n142 3328.24
R2767 dvdd.n216 dvdd.n140 3328.24
R2768 dvdd.n236 dvdd.n140 3328.24
R2769 dvdd.n562 dvdd.n557 2822.48
R2770 dvdd.n560 dvdd.n559 2822.48
R2771 dvdd.n596 dvdd.n263 2442.35
R2772 dvdd.n599 dvdd.n262 2442.35
R2773 dvdd.n569 dvdd.n554 2442.35
R2774 dvdd.n576 dvdd.n519 2442.35
R2775 dvdd.n584 dvdd.n583 2442.35
R2776 dvdd.n581 dvdd.n274 2442.35
R2777 dvdd.n44 dvdd.n43 2442.35
R2778 dvdd.n41 dvdd.n39 2442.35
R2779 dvdd.n32 dvdd.n31 2442.35
R2780 dvdd.n29 dvdd.n27 2442.35
R2781 dvdd.n20 dvdd.n19 2442.35
R2782 dvdd.n17 dvdd.n15 2442.35
R2783 dvdd.n8 dvdd.n7 2442.35
R2784 dvdd.n5 dvdd.n3 2442.35
R2785 dvdd.n194 dvdd.n122 1736.47
R2786 dvdd.n175 dvdd.n155 1736.47
R2787 dvdd.n225 dvdd.n160 1736.47
R2788 dvdd.n254 dvdd.n124 1736.47
R2789 dvdd.n602 dvdd.n106 1736.47
R2790 dvdd.n86 dvdd.n80 1736.47
R2791 dvdd.n617 dvdd.n104 1736.47
R2792 dvdd.n649 dvdd.n78 1736.47
R2793 dvdd.n574 dvdd.n522 1563.53
R2794 dvdd.n569 dvdd.n522 1563.53
R2795 dvdd.n576 dvdd.n520 1563.53
R2796 dvdd.n567 dvdd.n520 1563.53
R2797 dvdd.n268 dvdd.n266 1068.61
R2798 dvdd.n591 dvdd.n590 1068.61
R2799 dvdd.n201 dvdd.n200 878.823
R2800 dvdd.n200 dvdd.n170 878.823
R2801 dvdd.n173 dvdd.n163 878.823
R2802 dvdd.n174 dvdd.n173 878.823
R2803 dvdd.n202 dvdd.n169 878.823
R2804 dvdd.n202 dvdd.n201 878.823
R2805 dvdd.n145 dvdd.n123 878.823
R2806 dvdd.n244 dvdd.n123 878.823
R2807 dvdd.n209 dvdd.n208 878.823
R2808 dvdd.n208 dvdd.n163 878.823
R2809 dvdd.n168 dvdd.n132 878.823
R2810 dvdd.n169 dvdd.n168 878.823
R2811 dvdd.n236 dvdd.n234 878.823
R2812 dvdd.n234 dvdd.n147 878.823
R2813 dvdd.n214 dvdd.n213 878.823
R2814 dvdd.n214 dvdd.n153 878.823
R2815 dvdd.n210 dvdd.n153 878.823
R2816 dvdd.n210 dvdd.n209 878.823
R2817 dvdd.n216 dvdd.n152 878.823
R2818 dvdd.n227 dvdd.n152 878.823
R2819 dvdd.n228 dvdd.n227 878.823
R2820 dvdd.n228 dvdd.n132 878.823
R2821 dvdd.n147 dvdd.n130 878.823
R2822 dvdd.n243 dvdd.n130 878.823
R2823 dvdd.n243 dvdd.n131 878.823
R2824 dvdd.n182 dvdd.n131 878.823
R2825 dvdd.n244 dvdd.n121 878.823
R2826 dvdd.n121 dvdd.n118 878.823
R2827 dvdd.n256 dvdd.n118 878.823
R2828 dvdd.n256 dvdd.n119 878.823
R2829 dvdd.n182 dvdd.n180 878.823
R2830 dvdd.n191 dvdd.n180 878.823
R2831 dvdd.n192 dvdd.n191 878.823
R2832 dvdd.n193 dvdd.n192 878.823
R2833 dvdd.n122 dvdd.n119 878.823
R2834 dvdd.n175 dvdd.n174 878.823
R2835 dvdd.n237 dvdd.n142 878.823
R2836 dvdd.n237 dvdd.n236 878.823
R2837 dvdd.n217 dvdd.n141 878.823
R2838 dvdd.n217 dvdd.n216 878.823
R2839 dvdd.n254 dvdd.n125 878.823
R2840 dvdd.n125 dvdd.n120 878.823
R2841 dvdd.n145 dvdd.n120 878.823
R2842 dvdd.n213 dvdd.n160 878.823
R2843 dvdd.n65 dvdd.n54 878.823
R2844 dvdd.n65 dvdd.n61 878.823
R2845 dvdd.n608 dvdd.n109 878.823
R2846 dvdd.n608 dvdd.n607 878.823
R2847 dvdd.n611 dvdd.n111 878.823
R2848 dvdd.n611 dvdd.n94 878.823
R2849 dvdd.n95 dvdd.n60 878.823
R2850 dvdd.n96 dvdd.n95 878.823
R2851 dvdd.n542 dvdd.n61 878.823
R2852 dvdd.n543 dvdd.n542 878.823
R2853 dvdd.n607 dvdd.n606 878.823
R2854 dvdd.n606 dvdd.n115 878.823
R2855 dvdd.n532 dvdd.n94 878.823
R2856 dvdd.n533 dvdd.n532 878.823
R2857 dvdd.n526 dvdd.n96 878.823
R2858 dvdd.n527 dvdd.n526 878.823
R2859 dvdd.n544 dvdd.n543 878.823
R2860 dvdd.n545 dvdd.n544 878.823
R2861 dvdd.n602 dvdd.n115 878.823
R2862 dvdd.n535 dvdd.n533 878.823
R2863 dvdd.n535 dvdd.n534 878.823
R2864 dvdd.n529 dvdd.n527 878.823
R2865 dvdd.n529 dvdd.n528 878.823
R2866 dvdd.n547 dvdd.n545 878.823
R2867 dvdd.n547 dvdd.n546 878.823
R2868 dvdd.n86 dvdd.n85 878.823
R2869 dvdd.n636 dvdd.n632 878.823
R2870 dvdd.n636 dvdd.n635 878.823
R2871 dvdd.n635 dvdd.n634 878.823
R2872 dvdd.n634 dvdd.n633 878.823
R2873 dvdd.n644 dvdd.n83 878.823
R2874 dvdd.n644 dvdd.n643 878.823
R2875 dvdd.n643 dvdd.n642 878.823
R2876 dvdd.n642 dvdd.n85 878.823
R2877 dvdd.n62 dvdd.n53 878.823
R2878 dvdd.n62 dvdd.n60 878.823
R2879 dvdd.n110 dvdd.n101 878.823
R2880 dvdd.n111 dvdd.n110 878.823
R2881 dvdd.n109 dvdd.n104 878.823
R2882 dvdd.n75 dvdd.n74 878.823
R2883 dvdd.n75 dvdd.n69 878.823
R2884 dvdd.n631 dvdd.n69 878.823
R2885 dvdd.n632 dvdd.n631 878.823
R2886 dvdd.n83 dvdd.n78 878.823
R2887 dvdd.n524 dvdd.n522 878.823
R2888 dvdd.n524 dvdd.n520 878.823
R2889 dvdd.n226 dvdd.n153 857.648
R2890 dvdd.n227 dvdd.n226 857.648
R2891 dvdd.n147 dvdd.n146 857.648
R2892 dvdd.n146 dvdd.n145 857.648
R2893 dvdd.n209 dvdd.n158 857.648
R2894 dvdd.n158 dvdd.n132 857.648
R2895 dvdd.n245 dvdd.n243 857.648
R2896 dvdd.n245 dvdd.n244 857.648
R2897 dvdd.n163 dvdd.n157 857.648
R2898 dvdd.n169 dvdd.n157 857.648
R2899 dvdd.n183 dvdd.n182 857.648
R2900 dvdd.n183 dvdd.n118 857.648
R2901 dvdd.n174 dvdd.n156 857.648
R2902 dvdd.n201 dvdd.n156 857.648
R2903 dvdd.n191 dvdd.n190 857.648
R2904 dvdd.n190 dvdd.n119 857.648
R2905 dvdd.n170 dvdd.n155 857.648
R2906 dvdd.n194 dvdd.n193 857.648
R2907 dvdd.n225 dvdd.n141 857.648
R2908 dvdd.n142 dvdd.n124 857.648
R2909 dvdd.n213 dvdd.n159 857.648
R2910 dvdd.n216 dvdd.n159 857.648
R2911 dvdd.n236 dvdd.n235 857.648
R2912 dvdd.n235 dvdd.n125 857.648
R2913 dvdd.n534 dvdd.n106 857.648
R2914 dvdd.n633 dvdd.n80 857.648
R2915 dvdd.n115 dvdd.n107 857.648
R2916 dvdd.n533 dvdd.n107 857.648
R2917 dvdd.n635 dvdd.n81 857.648
R2918 dvdd.n85 dvdd.n81 857.648
R2919 dvdd.n607 dvdd.n108 857.648
R2920 dvdd.n108 dvdd.n94 857.648
R2921 dvdd.n632 dvdd.n82 857.648
R2922 dvdd.n643 dvdd.n82 857.648
R2923 dvdd.n617 dvdd.n101 857.648
R2924 dvdd.n649 dvdd.n74 857.648
R2925 dvdd.n616 dvdd.n109 857.648
R2926 dvdd.n616 dvdd.n111 857.648
R2927 dvdd.n648 dvdd.n69 857.648
R2928 dvdd.n648 dvdd.n83 857.648
R2929 dvdd.t16 dvdd.n97 741.205
R2930 dvdd.t16 dvdd.n55 741.205
R2931 dvdd.t13 dvdd.n55 741.205
R2932 dvdd.t13 dvdd.n56 741.205
R2933 dvdd.t18 dvdd.n56 741.205
R2934 dvdd.t18 dvdd.n70 741.205
R2935 dvdd.t2 dvdd.n521 659.64
R2936 dvdd.t118 dvdd.n521 659.64
R2937 dvdd.n552 dvdd.n551 656.188
R2938 dvdd.n551 dvdd.n550 656.188
R2939 dvdd.n538 dvdd.n537 656.188
R2940 dvdd.n539 dvdd.n538 656.188
R2941 dvdd.n540 dvdd.n539 656.188
R2942 dvdd.n541 dvdd.n540 656.188
R2943 dvdd.n541 dvdd.n89 656.188
R2944 dvdd.n638 dvdd.n89 656.188
R2945 dvdd.n623 dvdd.n93 656.188
R2946 dvdd.n624 dvdd.n623 656.188
R2947 dvdd.n625 dvdd.n624 656.188
R2948 dvdd.n626 dvdd.n625 656.188
R2949 dvdd.n627 dvdd.n626 656.188
R2950 dvdd.n629 dvdd.n627 656.188
R2951 dvdd.n614 dvdd.n613 656.188
R2952 dvdd.n613 dvdd.n64 656.188
R2953 dvdd.n657 dvdd.n64 656.188
R2954 dvdd.n657 dvdd.n656 656.188
R2955 dvdd.n656 dvdd.n655 656.188
R2956 dvdd.n655 dvdd.n68 656.188
R2957 dvdd.n563 dvdd.n556 545.13
R2958 dvdd.n556 dvdd.n275 545.13
R2959 dvdd.n575 dvdd.n519 535.419
R2960 dvdd.n568 dvdd.n554 535.419
R2961 dvdd.n274 dvdd.n272 535.419
R2962 dvdd.n583 dvdd.n582 535.419
R2963 dvdd.n39 dvdd.n38 535.419
R2964 dvdd.n43 dvdd.n42 535.419
R2965 dvdd.n27 dvdd.n26 535.419
R2966 dvdd.n31 dvdd.n30 535.419
R2967 dvdd.n15 dvdd.n14 535.419
R2968 dvdd.n19 dvdd.n18 535.419
R2969 dvdd.n3 dvdd.n2 535.419
R2970 dvdd.n7 dvdd.n6 535.419
R2971 dvdd.n553 dvdd.n552 436.104
R2972 dvdd.n240 dvdd.n143 355.012
R2973 dvdd.n240 dvdd.n239 355.012
R2974 dvdd.n220 dvdd.n219 355.012
R2975 dvdd.n219 dvdd.n144 355.012
R2976 dvdd.n231 dvdd.n230 355.012
R2977 dvdd.n232 dvdd.n231 355.012
R2978 dvdd.n151 dvdd.n133 355.012
R2979 dvdd.n133 dvdd.n129 355.012
R2980 dvdd.n204 dvdd.n166 355.012
R2981 dvdd.n185 dvdd.n166 355.012
R2982 dvdd.n187 dvdd.n167 355.012
R2983 dvdd.n188 dvdd.n187 355.012
R2984 dvdd.n198 dvdd.n197 355.012
R2985 dvdd.n197 dvdd.n196 355.012
R2986 dvdd.n594 dvdd.n593 348.613
R2987 dvdd.n593 dvdd.n265 348.613
R2988 dvdd.n559 dvdd.n558 318.108
R2989 dvdd.n562 dvdd.n561 318.108
R2990 dvdd.n565 dvdd.n563 295.529
R2991 dvdd.n578 dvdd.n275 295.529
R2992 dvdd.t6 dvdd.n134 271.635
R2993 dvdd.t6 dvdd.n135 271.635
R2994 dvdd.n40 dvdd.n36 260.519
R2995 dvdd.n28 dvdd.n24 260.519
R2996 dvdd.n16 dvdd.n12 260.519
R2997 dvdd.n4 dvdd.n0 260.519
R2998 dvdd.n600 dvdd.n261 260.329
R2999 dvdd.n601 dvdd.n600 243.018
R3000 dvdd.n594 dvdd.n261 229.702
R3001 dvdd.n422 dvdd.t25 229.419
R3002 dvdd.n477 dvdd.t19 229.419
R3003 dvdd.n48 dvdd.t14 229.419
R3004 dvdd.n508 dvdd.t3 229.212
R3005 dvdd.n505 dvdd.t11 229.212
R3006 dvdd.n507 dvdd.t115 229.179
R3007 dvdd.n417 dvdd.t12 229.076
R3008 dvdd.n47 dvdd.t5 228.484
R3009 dvdd.n35 dvdd.t22 228.484
R3010 dvdd.n23 dvdd.t117 228.484
R3011 dvdd.n11 dvdd.t1 228.484
R3012 dvdd.n422 dvdd.t17 228.215
R3013 dvdd.n298 dvdd.t74 228.215
R3014 dvdd.n419 dvdd.t7 228.215
R3015 dvdd.n418 dvdd.t8 228.215
R3016 dvdd.n417 dvdd.t9 228.215
R3017 dvdd.n294 dvdd.t83 228.215
R3018 dvdd.n495 dvdd.t98 228.215
R3019 dvdd.n398 dvdd.t54 228.215
R3020 dvdd.n283 dvdd.t40 228.215
R3021 dvdd.n510 dvdd.t50 228.215
R3022 dvdd.n514 dvdd.t51 228.215
R3023 dvdd.n517 dvdd.t119 228.215
R3024 dvdd.n278 dvdd.t67 228.215
R3025 dvdd.n452 dvdd.t48 228.215
R3026 dvdd.n454 dvdd.t47 228.215
R3027 dvdd.n450 dvdd.t44 228.215
R3028 dvdd.n448 dvdd.t45 228.215
R3029 dvdd.n446 dvdd.t94 228.215
R3030 dvdd.n444 dvdd.t95 228.215
R3031 dvdd.n435 dvdd.t76 228.215
R3032 dvdd.n433 dvdd.t77 228.215
R3033 dvdd.n477 dvdd.t120 228.215
R3034 dvdd.n48 dvdd.t20 228.215
R3035 dvdd.n431 dvdd.t80 228.215
R3036 dvdd.n428 dvdd.t79 228.215
R3037 dvdd.n436 dvdd.t89 228.215
R3038 dvdd.n437 dvdd.t88 228.215
R3039 dvdd.n455 dvdd.t68 228.215
R3040 dvdd.n281 dvdd.t41 228.215
R3041 dvdd.n383 dvdd.t107 228.215
R3042 dvdd.n319 dvdd.t106 228.215
R3043 dvdd.n318 dvdd.t103 228.215
R3044 dvdd.n313 dvdd.t37 228.215
R3045 dvdd.n311 dvdd.t38 228.215
R3046 dvdd.n309 dvdd.t34 228.215
R3047 dvdd.n307 dvdd.t35 228.215
R3048 dvdd.n305 dvdd.t31 228.215
R3049 dvdd.n303 dvdd.t32 228.215
R3050 dvdd.n301 dvdd.t100 228.215
R3051 dvdd.n351 dvdd.t61 228.215
R3052 dvdd.n344 dvdd.t85 228.215
R3053 dvdd.n340 dvdd.t91 228.215
R3054 dvdd.n336 dvdd.t109 228.215
R3055 dvdd.n332 dvdd.t64 228.215
R3056 dvdd.n323 dvdd.t27 228.215
R3057 dvdd.n321 dvdd.t28 228.215
R3058 dvdd.n329 dvdd.t70 228.215
R3059 dvdd.n324 dvdd.t71 228.215
R3060 dvdd.n326 dvdd.t65 228.215
R3061 dvdd.n334 dvdd.t110 228.215
R3062 dvdd.n338 dvdd.t92 228.215
R3063 dvdd.n342 dvdd.t86 228.215
R3064 dvdd.n346 dvdd.t62 228.215
R3065 dvdd.n348 dvdd.t112 228.215
R3066 dvdd.n355 dvdd.t113 228.215
R3067 dvdd.n299 dvdd.t101 228.215
R3068 dvdd.n397 dvdd.t104 228.215
R3069 dvdd.n385 dvdd.t57 228.215
R3070 dvdd.n284 dvdd.t58 228.215
R3071 dvdd.n286 dvdd.t55 228.215
R3072 dvdd.n291 dvdd.t97 228.215
R3073 dvdd.n292 dvdd.t82 228.215
R3074 dvdd.n295 dvdd.t73 228.215
R3075 dvdd.n597 dvdd.n596 214.912
R3076 dvdd.n599 dvdd.n598 214.912
R3077 dvdd.n177 dvdd.n176 185.225
R3078 dvdd.n224 dvdd.n223 185.225
R3079 dvdd.n549 dvdd.n87 185.225
R3080 dvdd.n40 dvdd.n37 176.139
R3081 dvdd.n28 dvdd.n25 176.139
R3082 dvdd.n16 dvdd.n13 176.139
R3083 dvdd.n4 dvdd.n1 176.139
R3084 dvdd.n603 dvdd.n601 167.906
R3085 dvdd.n580 dvdd.n265 160.376
R3086 dvdd.n580 dvdd.n579 160.376
R3087 dvdd.t81 dvdd.n489 120.174
R3088 dvdd.n490 dvdd.t81 120.174
R3089 dvdd.n493 dvdd.t96 120.174
R3090 dvdd.t96 dvdd.n289 120.174
R3091 dvdd.n462 dvdd.t46 120.174
R3092 dvdd.t46 dvdd.n461 120.174
R3093 dvdd.t42 dvdd.n465 120.174
R3094 dvdd.n466 dvdd.t42 120.174
R3095 dvdd.t93 dvdd.n469 120.174
R3096 dvdd.n470 dvdd.t93 120.174
R3097 dvdd.t75 dvdd.n473 120.174
R3098 dvdd.n474 dvdd.t75 120.174
R3099 dvdd.t56 dvdd.n285 120.174
R3100 dvdd.n388 dvdd.t56 120.174
R3101 dvdd.t105 dvdd.n391 120.174
R3102 dvdd.n392 dvdd.t105 120.174
R3103 dvdd.t33 dvdd.n406 120.174
R3104 dvdd.n407 dvdd.t33 120.174
R3105 dvdd.t29 dvdd.n410 120.174
R3106 dvdd.n411 dvdd.t29 120.174
R3107 dvdd.t99 dvdd.n414 120.174
R3108 dvdd.n415 dvdd.t99 120.174
R3109 dvdd.n352 dvdd.t59 120.174
R3110 dvdd.t59 dvdd.n347 120.174
R3111 dvdd.t84 dvdd.n362 120.174
R3112 dvdd.n363 dvdd.t84 120.174
R3113 dvdd.t90 dvdd.n366 120.174
R3114 dvdd.n367 dvdd.t90 120.174
R3115 dvdd.t108 dvdd.n370 120.174
R3116 dvdd.n371 dvdd.t108 120.174
R3117 dvdd.t63 dvdd.n374 120.174
R3118 dvdd.n375 dvdd.t63 120.174
R3119 dvdd.t69 dvdd.n325 120.174
R3120 dvdd.n328 dvdd.t69 120.174
R3121 dvdd.n403 dvdd.t36 120.174
R3122 dvdd.t36 dvdd.n402 120.174
R3123 dvdd.t102 dvdd.n315 120.174
R3124 dvdd.n395 dvdd.t102 120.174
R3125 dvdd.n499 dvdd.t52 120.174
R3126 dvdd.t52 dvdd.n498 120.174
R3127 dvdd.n46 dvdd.n36 118.127
R3128 dvdd.n34 dvdd.n24 118.127
R3129 dvdd.n22 dvdd.n12 118.127
R3130 dvdd.n10 dvdd.n0 118.127
R3131 dvdd.t53 dvdd.n105 103.335
R3132 dvdd.t53 dvdd.n97 103.335
R3133 dvdd.t43 dvdd.n70 103.335
R3134 dvdd.t43 dvdd.n79 103.335
R3135 dvdd.n610 dvdd.n112 100.141
R3136 dvdd.n610 dvdd.n609 100.141
R3137 dvdd.n609 dvdd.n114 100.141
R3138 dvdd.n605 dvdd.n604 100.141
R3139 dvdd.n604 dvdd.n603 100.141
R3140 dvdd.n536 dvdd.n270 98.7449
R3141 dvdd.n650 dvdd.n77 96.5745
R3142 dvdd.n222 dvdd.n215 93.7417
R3143 dvdd.n215 dvdd.n212 93.7417
R3144 dvdd.n212 dvdd.n211 93.7417
R3145 dvdd.n211 dvdd.n162 93.7417
R3146 dvdd.n207 dvdd.n162 93.7417
R3147 dvdd.n207 dvdd.n206 93.7417
R3148 dvdd.n206 dvdd.n164 93.7417
R3149 dvdd.n172 dvdd.n164 93.7417
R3150 dvdd.n176 dvdd.n172 93.7417
R3151 dvdd.n239 dvdd.n238 93.7417
R3152 dvdd.n238 dvdd.n144 93.7417
R3153 dvdd.n223 dvdd.n222 93.7417
R3154 dvdd.n218 dvdd.n143 93.7417
R3155 dvdd.n220 dvdd.n218 93.7417
R3156 dvdd.n220 dvdd.n149 93.7417
R3157 dvdd.n230 dvdd.n149 93.7417
R3158 dvdd.n233 dvdd.n144 93.7417
R3159 dvdd.n233 dvdd.n232 93.7417
R3160 dvdd.n232 dvdd.n148 93.7417
R3161 dvdd.n148 dvdd.n129 93.7417
R3162 dvdd.n230 dvdd.n229 93.7417
R3163 dvdd.n229 dvdd.n151 93.7417
R3164 dvdd.n165 dvdd.n151 93.7417
R3165 dvdd.n204 dvdd.n165 93.7417
R3166 dvdd.n181 dvdd.n129 93.7417
R3167 dvdd.n185 dvdd.n181 93.7417
R3168 dvdd.n186 dvdd.n185 93.7417
R3169 dvdd.n188 dvdd.n186 93.7417
R3170 dvdd.n204 dvdd.n203 93.7417
R3171 dvdd.n203 dvdd.n167 93.7417
R3172 dvdd.n199 dvdd.n167 93.7417
R3173 dvdd.n199 dvdd.n198 93.7417
R3174 dvdd.n188 dvdd.n178 93.7417
R3175 dvdd.n196 dvdd.n178 93.7417
R3176 dvdd.n651 dvdd.n76 93.7417
R3177 dvdd.n76 dvdd.n68 93.7417
R3178 dvdd.n66 dvdd.n52 93.7417
R3179 dvdd.n656 dvdd.n66 93.7417
R3180 dvdd.n614 dvdd.n612 93.7417
R3181 dvdd.n612 dvdd.n93 93.7417
R3182 dvdd.n91 dvdd.n64 93.7417
R3183 dvdd.n624 dvdd.n91 93.7417
R3184 dvdd.n656 dvdd.n67 93.7417
R3185 dvdd.n626 dvdd.n67 93.7417
R3186 dvdd.n531 dvdd.n93 93.7417
R3187 dvdd.n537 dvdd.n531 93.7417
R3188 dvdd.n537 dvdd.n536 93.7417
R3189 dvdd.n624 dvdd.n92 93.7417
R3190 dvdd.n539 dvdd.n92 93.7417
R3191 dvdd.n539 dvdd.n530 93.7417
R3192 dvdd.n530 dvdd.n271 93.7417
R3193 dvdd.n626 dvdd.n90 93.7417
R3194 dvdd.n541 dvdd.n90 93.7417
R3195 dvdd.n548 dvdd.n541 93.7417
R3196 dvdd.n552 dvdd.n548 93.7417
R3197 dvdd.n638 dvdd.n88 93.7417
R3198 dvdd.n550 dvdd.n88 93.7417
R3199 dvdd.n641 dvdd.n84 93.7417
R3200 dvdd.n641 dvdd.n640 93.7417
R3201 dvdd.n640 dvdd.n87 93.7417
R3202 dvdd.n630 dvdd.n68 93.7417
R3203 dvdd.n630 dvdd.n629 93.7417
R3204 dvdd.n637 dvdd.n629 93.7417
R3205 dvdd.n638 dvdd.n637 93.7417
R3206 dvdd.n63 dvdd.n51 93.7417
R3207 dvdd.n64 dvdd.n63 93.7417
R3208 dvdd.n646 dvdd.n77 93.7417
R3209 dvdd.n646 dvdd.n645 93.7417
R3210 dvdd.n645 dvdd.n84 93.7417
R3211 dvdd.n619 dvdd.n102 93.7417
R3212 dvdd.n614 dvdd.n102 93.7417
R3213 dvdd.n112 dvdd.n103 93.7417
R3214 dvdd.n605 dvdd.n258 93.7417
R3215 dvdd.n572 dvdd.n525 93.7417
R3216 dvdd.n555 dvdd.n525 93.7417
R3217 dvdd.n253 dvdd.n126 91.6685
R3218 dvdd.n195 dvdd.n179 91.6685
R3219 dvdd.n224 dvdd.n143 91.4829
R3220 dvdd.n239 dvdd.n126 91.4829
R3221 dvdd.n222 dvdd.n221 91.4829
R3222 dvdd.n221 dvdd.n220 91.4829
R3223 dvdd.n144 dvdd.n127 91.4829
R3224 dvdd.n212 dvdd.n150 91.4829
R3225 dvdd.n230 dvdd.n150 91.4829
R3226 dvdd.n232 dvdd.n128 91.4829
R3227 dvdd.n162 dvdd.n161 91.4829
R3228 dvdd.n161 dvdd.n151 91.4829
R3229 dvdd.n246 dvdd.n129 91.4829
R3230 dvdd.n206 dvdd.n205 91.4829
R3231 dvdd.n205 dvdd.n204 91.4829
R3232 dvdd.n185 dvdd.n184 91.4829
R3233 dvdd.n172 dvdd.n171 91.4829
R3234 dvdd.n171 dvdd.n167 91.4829
R3235 dvdd.n189 dvdd.n188 91.4829
R3236 dvdd.n198 dvdd.n177 91.4829
R3237 dvdd.n196 dvdd.n195 91.4829
R3238 dvdd.n550 dvdd.n549 91.4829
R3239 dvdd.n537 dvdd.n259 91.4829
R3240 dvdd.n639 dvdd.n638 91.4829
R3241 dvdd.n640 dvdd.n639 91.4829
R3242 dvdd.n113 dvdd.n93 91.4829
R3243 dvdd.n629 dvdd.n628 91.4829
R3244 dvdd.n628 dvdd.n84 91.4829
R3245 dvdd.n615 dvdd.n614 91.4829
R3246 dvdd.n647 dvdd.n68 91.4829
R3247 dvdd.n647 dvdd.n646 91.4829
R3248 dvdd.n252 dvdd.n127 85.0829
R3249 dvdd.n250 dvdd.n128 85.0829
R3250 dvdd.n248 dvdd.n246 85.0829
R3251 dvdd.n184 dvdd.n116 85.0829
R3252 dvdd.n189 dvdd.n117 85.0829
R3253 dvdd.n604 dvdd.n259 85.0829
R3254 dvdd.n114 dvdd.n113 85.0829
R3255 dvdd.n615 dvdd.n610 85.0829
R3256 dvdd.n386 dvdd.t24 84.9815
R3257 dvdd.t60 dvdd.n154 69.9975
R3258 dvdd.t60 dvdd.n134 69.9975
R3259 dvdd.n135 dvdd.t30 69.9975
R3260 dvdd.n255 dvdd.t30 69.9975
R3261 dvdd.n579 dvdd.n578 44.796
R3262 dvdd.n45 dvdd.n37 44.2181
R3263 dvdd.n33 dvdd.n25 44.2181
R3264 dvdd.n21 dvdd.n13 44.2181
R3265 dvdd.n9 dvdd.n1 44.2181
R3266 dvdd.n565 dvdd.n564 38.4243
R3267 dvdd.n225 dvdd.n224 37.0005
R3268 dvdd.t60 dvdd.n225 37.0005
R3269 dvdd.n126 dvdd.n124 37.0005
R3270 dvdd.n124 dvdd.t30 37.0005
R3271 dvdd.n221 dvdd.n159 37.0005
R3272 dvdd.t60 dvdd.n159 37.0005
R3273 dvdd.n235 dvdd.n127 37.0005
R3274 dvdd.n235 dvdd.t30 37.0005
R3275 dvdd.n226 dvdd.n150 37.0005
R3276 dvdd.n226 dvdd.t60 37.0005
R3277 dvdd.n146 dvdd.n128 37.0005
R3278 dvdd.n146 dvdd.t30 37.0005
R3279 dvdd.n161 dvdd.n158 37.0005
R3280 dvdd.t60 dvdd.n158 37.0005
R3281 dvdd.n246 dvdd.n245 37.0005
R3282 dvdd.n245 dvdd.t30 37.0005
R3283 dvdd.n205 dvdd.n157 37.0005
R3284 dvdd.t60 dvdd.n157 37.0005
R3285 dvdd.n184 dvdd.n183 37.0005
R3286 dvdd.n183 dvdd.t30 37.0005
R3287 dvdd.n171 dvdd.n156 37.0005
R3288 dvdd.t60 dvdd.n156 37.0005
R3289 dvdd.n190 dvdd.n189 37.0005
R3290 dvdd.n190 dvdd.t30 37.0005
R3291 dvdd.n195 dvdd.n194 37.0005
R3292 dvdd.n194 dvdd.t30 37.0005
R3293 dvdd.n177 dvdd.n155 37.0005
R3294 dvdd.t60 dvdd.n155 37.0005
R3295 dvdd.n262 dvdd.n260 37.0005
R3296 dvdd.n113 dvdd.n108 37.0005
R3297 dvdd.t53 dvdd.n108 37.0005
R3298 dvdd.n259 dvdd.n107 37.0005
R3299 dvdd.t53 dvdd.n107 37.0005
R3300 dvdd.n628 dvdd.n82 37.0005
R3301 dvdd.t43 dvdd.n82 37.0005
R3302 dvdd.n639 dvdd.n81 37.0005
R3303 dvdd.t43 dvdd.n81 37.0005
R3304 dvdd.n549 dvdd.n80 37.0005
R3305 dvdd.t43 dvdd.n80 37.0005
R3306 dvdd.n269 dvdd.n106 37.0005
R3307 dvdd.t53 dvdd.n106 37.0005
R3308 dvdd.n616 dvdd.n615 37.0005
R3309 dvdd.t53 dvdd.n616 37.0005
R3310 dvdd.n648 dvdd.n647 37.0005
R3311 dvdd.t43 dvdd.n648 37.0005
R3312 dvdd.n618 dvdd.n617 37.0005
R3313 dvdd.n617 dvdd.t53 37.0005
R3314 dvdd.n650 dvdd.n649 37.0005
R3315 dvdd.n649 dvdd.t43 37.0005
R3316 dvdd.n263 dvdd.n261 37.0005
R3317 dvdd.n597 dvdd.n262 33.2417
R3318 dvdd.n598 dvdd.n263 33.2417
R3319 dvdd.n564 dvdd.n553 31.2476
R3320 dvdd.n176 dvdd.n175 30.8338
R3321 dvdd.n175 dvdd.n154 30.8338
R3322 dvdd.n173 dvdd.n164 30.8338
R3323 dvdd.n173 dvdd.n154 30.8338
R3324 dvdd.n208 dvdd.n207 30.8338
R3325 dvdd.n208 dvdd.n154 30.8338
R3326 dvdd.n211 dvdd.n210 30.8338
R3327 dvdd.n210 dvdd.n154 30.8338
R3328 dvdd.n215 dvdd.n214 30.8338
R3329 dvdd.n214 dvdd.n154 30.8338
R3330 dvdd.n238 dvdd.n237 30.8338
R3331 dvdd.n237 dvdd.n135 30.8338
R3332 dvdd.n223 dvdd.n160 30.8338
R3333 dvdd.n160 dvdd.n154 30.8338
R3334 dvdd.n218 dvdd.n217 30.8338
R3335 dvdd.n217 dvdd.n134 30.8338
R3336 dvdd.n152 dvdd.n149 30.8338
R3337 dvdd.n152 dvdd.n134 30.8338
R3338 dvdd.n234 dvdd.n233 30.8338
R3339 dvdd.n234 dvdd.n135 30.8338
R3340 dvdd.n148 dvdd.n130 30.8338
R3341 dvdd.n135 dvdd.n130 30.8338
R3342 dvdd.n229 dvdd.n228 30.8338
R3343 dvdd.n228 dvdd.n134 30.8338
R3344 dvdd.n168 dvdd.n165 30.8338
R3345 dvdd.n168 dvdd.n134 30.8338
R3346 dvdd.n181 dvdd.n131 30.8338
R3347 dvdd.n135 dvdd.n131 30.8338
R3348 dvdd.n186 dvdd.n180 30.8338
R3349 dvdd.n180 dvdd.n135 30.8338
R3350 dvdd.n203 dvdd.n202 30.8338
R3351 dvdd.n202 dvdd.n134 30.8338
R3352 dvdd.n200 dvdd.n199 30.8338
R3353 dvdd.n200 dvdd.n134 30.8338
R3354 dvdd.n192 dvdd.n178 30.8338
R3355 dvdd.n192 dvdd.n135 30.8338
R3356 dvdd.n254 dvdd.n253 30.8338
R3357 dvdd.n255 dvdd.n254 30.8338
R3358 dvdd.n251 dvdd.n120 30.8338
R3359 dvdd.n255 dvdd.n120 30.8338
R3360 dvdd.n249 dvdd.n123 30.8338
R3361 dvdd.n255 dvdd.n123 30.8338
R3362 dvdd.n247 dvdd.n121 30.8338
R3363 dvdd.n255 dvdd.n121 30.8338
R3364 dvdd.n257 dvdd.n256 30.8338
R3365 dvdd.n256 dvdd.n255 30.8338
R3366 dvdd.n179 dvdd.n122 30.8338
R3367 dvdd.n255 dvdd.n122 30.8338
R3368 dvdd.n634 dvdd.n88 30.8338
R3369 dvdd.n634 dvdd.n70 30.8338
R3370 dvdd.n548 dvdd.n547 30.8338
R3371 dvdd.n547 dvdd.n56 30.8338
R3372 dvdd.n530 dvdd.n529 30.8338
R3373 dvdd.n529 dvdd.n55 30.8338
R3374 dvdd.n66 dvdd.n65 30.8338
R3375 dvdd.n65 dvdd.n56 30.8338
R3376 dvdd.n542 dvdd.n67 30.8338
R3377 dvdd.n542 dvdd.n56 30.8338
R3378 dvdd.n95 dvdd.n91 30.8338
R3379 dvdd.n95 dvdd.n55 30.8338
R3380 dvdd.n612 dvdd.n611 30.8338
R3381 dvdd.n611 dvdd.n97 30.8338
R3382 dvdd.n642 dvdd.n641 30.8338
R3383 dvdd.n642 dvdd.n79 30.8338
R3384 dvdd.n637 dvdd.n636 30.8338
R3385 dvdd.n636 dvdd.n70 30.8338
R3386 dvdd.n544 dvdd.n90 30.8338
R3387 dvdd.n544 dvdd.n56 30.8338
R3388 dvdd.n526 dvdd.n92 30.8338
R3389 dvdd.n526 dvdd.n55 30.8338
R3390 dvdd.n532 dvdd.n531 30.8338
R3391 dvdd.n532 dvdd.n97 30.8338
R3392 dvdd.n536 dvdd.n535 30.8338
R3393 dvdd.n535 dvdd.n97 30.8338
R3394 dvdd.n87 dvdd.n86 30.8338
R3395 dvdd.n86 dvdd.n79 30.8338
R3396 dvdd.n63 dvdd.n62 30.8338
R3397 dvdd.n62 dvdd.n55 30.8338
R3398 dvdd.n76 dvdd.n75 30.8338
R3399 dvdd.n75 dvdd.n70 30.8338
R3400 dvdd.n631 dvdd.n630 30.8338
R3401 dvdd.n631 dvdd.n70 30.8338
R3402 dvdd.n78 dvdd.n77 30.8338
R3403 dvdd.n79 dvdd.n78 30.8338
R3404 dvdd.n645 dvdd.n644 30.8338
R3405 dvdd.n644 dvdd.n79 30.8338
R3406 dvdd.n110 dvdd.n102 30.8338
R3407 dvdd.n110 dvdd.n97 30.8338
R3408 dvdd.n603 dvdd.n602 30.8338
R3409 dvdd.n602 dvdd.n105 30.8338
R3410 dvdd.n606 dvdd.n605 30.8338
R3411 dvdd.n606 dvdd.n105 30.8338
R3412 dvdd.n609 dvdd.n608 30.8338
R3413 dvdd.n608 dvdd.n105 30.8338
R3414 dvdd.n112 dvdd.n104 30.8338
R3415 dvdd.n105 dvdd.n104 30.8338
R3416 dvdd.n268 dvdd.n264 30.8338
R3417 dvdd.n525 dvdd.n524 30.8338
R3418 dvdd.n524 dvdd.n521 30.8338
R3419 dvdd.n583 dvdd.n273 30.8338
R3420 dvdd.n519 dvdd.n273 30.8338
R3421 dvdd.n591 dvdd.n267 30.8338
R3422 dvdd.n274 dvdd.n267 30.8338
R3423 dvdd.n564 dvdd.n554 30.8338
R3424 dvdd.n43 dvdd.n37 30.8338
R3425 dvdd.n39 dvdd.n36 30.8338
R3426 dvdd.n31 dvdd.n25 30.8338
R3427 dvdd.n27 dvdd.n24 30.8338
R3428 dvdd.n19 dvdd.n13 30.8338
R3429 dvdd.n15 dvdd.n12 30.8338
R3430 dvdd.n7 dvdd.n1 30.8338
R3431 dvdd.n3 dvdd.n0 30.8338
R3432 dvdd.n588 dvdd.n270 30.0837
R3433 dvdd.n587 dvdd.n586 25.7304
R3434 dvdd.n620 dvdd.n619 20.3196
R3435 dvdd.n620 dvdd.n51 20.3196
R3436 dvdd.n660 dvdd.n52 20.3196
R3437 dvdd.n652 dvdd.n52 20.3196
R3438 dvdd.n652 dvdd.n651 20.3196
R3439 dvdd.n586 dvdd.n585 20.2401
R3440 dvdd.n573 dvdd.n523 20.2401
R3441 dvdd.n661 dvdd.n51 17.1488
R3442 dvdd.n600 dvdd.n599 16.8187
R3443 dvdd.n596 dvdd.n595 16.8187
R3444 dvdd.n581 dvdd.n580 16.8187
R3445 dvdd.n585 dvdd.n584 16.8187
R3446 dvdd.n574 dvdd.n573 16.8187
R3447 dvdd.n570 dvdd.n569 16.8187
R3448 dvdd.n569 dvdd.t118 16.8187
R3449 dvdd.n567 dvdd.n566 16.8187
R3450 dvdd.n577 dvdd.n576 16.8187
R3451 dvdd.n576 dvdd.t2 16.8187
R3452 dvdd.n41 dvdd.n40 16.8187
R3453 dvdd.n45 dvdd.n44 16.8187
R3454 dvdd.n29 dvdd.n28 16.8187
R3455 dvdd.n33 dvdd.n32 16.8187
R3456 dvdd.n17 dvdd.n16 16.8187
R3457 dvdd.n21 dvdd.n20 16.8187
R3458 dvdd.n5 dvdd.n4 16.8187
R3459 dvdd.n9 dvdd.n8 16.8187
R3460 dvdd.n570 dvdd.n553 15.4969
R3461 dvdd.n573 dvdd.n572 14.3924
R3462 dvdd.n575 dvdd.n574 13.0425
R3463 dvdd.n584 dvdd.n272 13.0425
R3464 dvdd.n582 dvdd.n581 13.0425
R3465 dvdd.n568 dvdd.n567 13.0425
R3466 dvdd.n44 dvdd.n38 13.0425
R3467 dvdd.n42 dvdd.n41 13.0425
R3468 dvdd.n32 dvdd.n26 13.0425
R3469 dvdd.n30 dvdd.n29 13.0425
R3470 dvdd.n20 dvdd.n14 13.0425
R3471 dvdd.n18 dvdd.n17 13.0425
R3472 dvdd.n8 dvdd.n2 13.0425
R3473 dvdd.n6 dvdd.n5 13.0425
R3474 dvdd.n572 dvdd.n571 12.4107
R3475 dvdd.t111 dvdd.n357 11.9724
R3476 dvdd.n358 dvdd.t111 11.9724
R3477 dvdd.t26 dvdd.n379 11.9724
R3478 dvdd.n380 dvdd.t26 11.9724
R3479 dvdd.n270 dvdd.n264 11.3275
R3480 dvdd.n560 dvdd.n556 10.8829
R3481 dvdd.n557 dvdd.n518 10.8829
R3482 dvdd.n588 dvdd.n587 10.7538
R3483 dvdd.n585 dvdd.n271 10.6563
R3484 dvdd.n566 dvdd.n555 9.69349
R3485 dvdd.n558 dvdd.n557 9.61977
R3486 dvdd.n561 dvdd.n560 9.61977
R3487 dvdd.n523 dvdd.n271 9.58426
R3488 dvdd.n563 dvdd.n562 8.81002
R3489 dvdd.n559 dvdd.n275 8.81002
R3490 dvdd.n579 dvdd.n273 8.64212
R3491 dvdd.n267 dvdd.n265 8.64212
R3492 dvdd.n577 dvdd.n518 8.13999
R3493 dvdd.n523 dvdd.n273 8.08984
R3494 dvdd.n586 dvdd.n267 8.08984
R3495 dvdd.n241 dvdd.n240 7.4005
R3496 dvdd.t6 dvdd.n241 7.4005
R3497 dvdd.n219 dvdd.n140 7.4005
R3498 dvdd.t6 dvdd.n140 7.4005
R3499 dvdd.n231 dvdd.n139 7.4005
R3500 dvdd.t6 dvdd.n139 7.4005
R3501 dvdd.n242 dvdd.n133 7.4005
R3502 dvdd.n242 dvdd.t6 7.4005
R3503 dvdd.n166 dvdd.n138 7.4005
R3504 dvdd.t6 dvdd.n138 7.4005
R3505 dvdd.n187 dvdd.n137 7.4005
R3506 dvdd.t6 dvdd.n137 7.4005
R3507 dvdd.n197 dvdd.n136 7.4005
R3508 dvdd.t6 dvdd.n136 7.4005
R3509 dvdd.n593 dvdd.n592 7.4005
R3510 dvdd.n589 dvdd.n588 7.4005
R3511 dvdd.n601 dvdd.n260 7.31014
R3512 dvdd.n270 dvdd.n269 7.31014
R3513 dvdd.n253 dvdd.n252 6.58619
R3514 dvdd.n252 dvdd.n251 6.58619
R3515 dvdd.n251 dvdd.n250 6.58619
R3516 dvdd.n250 dvdd.n249 6.58619
R3517 dvdd.n249 dvdd.n248 6.58619
R3518 dvdd.n248 dvdd.n247 6.58619
R3519 dvdd.n247 dvdd.n116 6.58619
R3520 dvdd.n257 dvdd.n117 6.58619
R3521 dvdd.n179 dvdd.n117 6.58619
R3522 dvdd.n258 dvdd.n114 6.4005
R3523 dvdd.n578 dvdd.n577 6.36768
R3524 dvdd.n258 dvdd.n257 6.1653
R3525 dvdd.n486 dvdd.t72 5.91616
R3526 dvdd.t72 dvdd.n485 5.91616
R3527 dvdd.t39 dvdd.n503 5.91616
R3528 dvdd.n504 dvdd.t39 5.91616
R3529 dvdd.n512 dvdd.t49 5.91616
R3530 dvdd.t49 dvdd.n276 5.91616
R3531 dvdd.n458 dvdd.t66 5.91616
R3532 dvdd.t66 dvdd.n457 5.91616
R3533 dvdd.t78 dvdd.n481 5.91616
R3534 dvdd.n482 dvdd.t78 5.91616
R3535 dvdd.t87 dvdd.n440 5.91616
R3536 dvdd.n441 dvdd.t87 5.91616
R3537 dvdd.n590 dvdd.n589 5.51167
R3538 dvdd.n592 dvdd.n266 5.51167
R3539 dvdd.n485 dvdd.n484 5.13093
R3540 dvdd.n595 dvdd.n264 5.07987
R3541 dvdd.n423 dvdd.n422 4.88319
R3542 dvdd.n478 dvdd.n477 4.88319
R3543 dvdd.n49 dvdd.n48 4.88319
R3544 dvdd.n441 dvdd.n438 4.42713
R3545 dvdd.n483 dvdd.n482 4.42713
R3546 dvdd.n457 dvdd.n279 4.42713
R3547 dvdd.n458 dvdd.n277 4.42713
R3548 dvdd.n512 dvdd.n511 4.42713
R3549 dvdd.n504 dvdd.n282 4.42713
R3550 dvdd.n503 dvdd.n502 4.42713
R3551 dvdd.n485 dvdd.n297 4.42713
R3552 dvdd.n487 dvdd.n486 4.42713
R3553 dvdd.n481 dvdd.n480 4.38659
R3554 dvdd.n481 dvdd.n430 4.37758
R3555 dvdd.n440 dvdd.n432 4.37758
R3556 dvdd.n440 dvdd.n439 4.36463
R3557 dvdd.n442 dvdd.n441 4.36463
R3558 dvdd.n482 dvdd.n429 4.36463
R3559 dvdd.n457 dvdd.n456 4.36463
R3560 dvdd.n459 dvdd.n458 4.36463
R3561 dvdd.n513 dvdd.n512 4.36463
R3562 dvdd.n503 dvdd.n280 4.36463
R3563 dvdd.n486 dvdd.n296 4.36463
R3564 dvdd.n627 dvdd.n73 3.77601
R3565 dvdd.t18 dvdd.n73 3.77601
R3566 dvdd.n625 dvdd.n59 3.77601
R3567 dvdd.t13 dvdd.n59 3.77601
R3568 dvdd.n623 dvdd.n622 3.77601
R3569 dvdd.n622 dvdd.t16 3.77601
R3570 dvdd.n538 dvdd.n99 3.77601
R3571 dvdd.t16 dvdd.n99 3.77601
R3572 dvdd.n540 dvdd.n58 3.77601
R3573 dvdd.t13 dvdd.n58 3.77601
R3574 dvdd.n89 dvdd.n72 3.77601
R3575 dvdd.t18 dvdd.n72 3.77601
R3576 dvdd.n551 dvdd.n71 3.77601
R3577 dvdd.t18 dvdd.n71 3.77601
R3578 dvdd.n613 dvdd.n100 3.77601
R3579 dvdd.t16 dvdd.n100 3.77601
R3580 dvdd.n658 dvdd.n657 3.77601
R3581 dvdd.t13 dvdd.n658 3.77601
R3582 dvdd.n655 dvdd.n654 3.77601
R3583 dvdd.n654 dvdd.t18 3.77601
R3584 dvdd.n621 dvdd.n620 3.77601
R3585 dvdd.t16 dvdd.n621 3.77601
R3586 dvdd.n660 dvdd.n659 3.77601
R3587 dvdd.n659 dvdd.t13 3.77601
R3588 dvdd.n653 dvdd.n652 3.77601
R3589 dvdd.t18 dvdd.n653 3.77601
R3590 dvdd.n571 dvdd.n57 3.77601
R3591 dvdd.t13 dvdd.n57 3.77601
R3592 dvdd.n587 dvdd.n98 3.77601
R3593 dvdd.t16 dvdd.n98 3.77601
R3594 dvdd.t118 dvdd.n568 3.68792
R3595 dvdd.n582 dvdd.t114 3.68792
R3596 dvdd.t114 dvdd.n272 3.68792
R3597 dvdd.t2 dvdd.n575 3.68792
R3598 dvdd.n42 dvdd.t4 3.68792
R3599 dvdd.t4 dvdd.n38 3.68792
R3600 dvdd.n30 dvdd.t21 3.68792
R3601 dvdd.t21 dvdd.n26 3.68792
R3602 dvdd.n18 dvdd.t116 3.68792
R3603 dvdd.t116 dvdd.n14 3.68792
R3604 dvdd.n6 dvdd.t0 3.68792
R3605 dvdd.t0 dvdd.n2 3.68792
R3606 dvdd.n566 dvdd.n565 3.26067
R3607 dvdd.n598 dvdd.t23 3.25677
R3608 dvdd.t23 dvdd.n597 3.25677
R3609 dvdd.n661 dvdd.n660 3.17136
R3610 dvdd.n509 dvdd.n508 3.10376
R3611 dvdd.n516 dvdd.n515 3.04126
R3612 dvdd.n618 dvdd.n103 2.83329
R3613 dvdd.n619 dvdd.n618 2.83329
R3614 dvdd.n651 dvdd.n650 2.83329
R3615 dvdd.n506 dvdd.n505 2.74778
R3616 dvdd.n665 dvdd.n664 2.66096
R3617 dvdd.n420 dvdd.n419 2.42664
R3618 dvdd.n380 dvdd.n322 2.25322
R3619 dvdd.n379 dvdd.n378 2.25322
R3620 dvdd.n359 dvdd.n358 2.25322
R3621 dvdd.n357 dvdd.n354 2.25322
R3622 dvdd.n358 dvdd.n349 2.19072
R3623 dvdd.n357 dvdd.n356 2.19072
R3624 dvdd.n381 dvdd.n380 2.188
R3625 dvdd.n379 dvdd.n320 2.188
R3626 dvdd.n390 dvdd.n389 2.02496
R3627 dvdd.n571 dvdd.n570 1.98223
R3628 dvdd.t10 dvdd.n266 1.88064
R3629 dvdd.n590 dvdd.t10 1.88064
R3630 dvdd.n595 dvdd.n594 1.67669
R3631 dvdd.n555 dvdd.n518 1.554
R3632 dvdd.n505 dvdd.n504 1.37822
R3633 dvdd.n518 dvdd 1.3042
R3634 dvdd.n561 dvdd.t15 1.2275
R3635 dvdd.n558 dvdd.t15 1.2275
R3636 dvdd dvdd.n517 1.19558
R3637 dvdd.n508 dvdd.n276 1.08474
R3638 dvdd.n516 dvdd.n276 1.08474
R3639 dvdd.n517 dvdd.n516 0.996712
R3640 dvdd.n298 dvdd.n296 0.891804
R3641 dvdd.n418 dvdd.n417 0.860794
R3642 dvdd.n419 dvdd.n418 0.84943
R3643 dvdd.n484 dvdd.n483 0.791063
R3644 dvdd.n424 dvdd 0.751032
R3645 dvdd.n461 dvdd.n452 0.734196
R3646 dvdd.n329 dvdd.n328 0.734196
R3647 dvdd.n352 dvdd.n351 0.734196
R3648 dvdd.n47 dvdd.n46 0.639894
R3649 dvdd.n35 dvdd.n34 0.639894
R3650 dvdd.n23 dvdd.n22 0.639894
R3651 dvdd.n11 dvdd.n10 0.639894
R3652 dvdd dvdd.n667 0.62021
R3653 dvdd.n327 dvdd.n322 0.620065
R3654 dvdd.n378 dvdd.n377 0.620065
R3655 dvdd.n360 dvdd.n359 0.620065
R3656 dvdd.n354 dvdd.n353 0.620065
R3657 dvdd.n502 dvdd.n501 0.620065
R3658 dvdd.n297 dvdd.n290 0.620065
R3659 dvdd.n488 dvdd.n487 0.620065
R3660 dvdd.n426 dvdd.n425 0.603761
R3661 dvdd.n664 dvdd.n663 0.549667
R3662 dvdd.n476 dvdd.n475 0.478761
R3663 dvdd.n386 dvdd.n282 0.478761
R3664 dvdd.n421 dvdd.n293 0.478761
R3665 dvdd.n426 dvdd.n296 0.478761
R3666 dvdd.n425 dvdd.n421 0.474712
R3667 dvdd.n460 dvdd.n459 0.470609
R3668 dvdd.n438 dvdd.n429 0.470609
R3669 dvdd.n439 dvdd.n434 0.470609
R3670 dvdd.n443 dvdd.n442 0.470609
R3671 dvdd.n456 dvdd.n453 0.470609
R3672 dvdd.n513 dvdd.n279 0.470609
R3673 dvdd.n515 dvdd.n277 0.470609
R3674 dvdd.n511 dvdd.n280 0.470609
R3675 dvdd.n666 dvdd.n665 0.464907
R3676 dvdd.n667 dvdd.n666 0.464907
R3677 dvdd.n384 dvdd.n287 0.429848
R3678 dvdd.n445 dvdd.n443 0.429848
R3679 dvdd.n472 dvdd.n471 0.429848
R3680 dvdd.n449 dvdd.n447 0.429848
R3681 dvdd.n468 dvdd.n467 0.429848
R3682 dvdd.n453 dvdd.n451 0.429848
R3683 dvdd.n464 dvdd.n463 0.429848
R3684 dvdd.n331 dvdd.n330 0.429848
R3685 dvdd.n377 dvdd.n376 0.429848
R3686 dvdd.n335 dvdd.n333 0.429848
R3687 dvdd.n373 dvdd.n372 0.429848
R3688 dvdd.n339 dvdd.n337 0.429848
R3689 dvdd.n369 dvdd.n368 0.429848
R3690 dvdd.n343 dvdd.n341 0.429848
R3691 dvdd.n365 dvdd.n364 0.429848
R3692 dvdd.n350 dvdd.n345 0.429848
R3693 dvdd.n361 dvdd.n360 0.429848
R3694 dvdd.n304 dvdd.n302 0.429848
R3695 dvdd.n413 dvdd.n412 0.429848
R3696 dvdd.n308 dvdd.n306 0.429848
R3697 dvdd.n409 dvdd.n408 0.429848
R3698 dvdd.n312 dvdd.n310 0.429848
R3699 dvdd.n405 dvdd.n404 0.429848
R3700 dvdd.n317 dvdd.n314 0.429848
R3701 dvdd.n396 dvdd.n316 0.429848
R3702 dvdd.n394 dvdd.n393 0.429848
R3703 dvdd.n497 dvdd.n496 0.429848
R3704 dvdd.n501 dvdd.n500 0.429848
R3705 dvdd.n494 dvdd.n290 0.429848
R3706 dvdd.n492 dvdd.n491 0.429848
R3707 dvdd.n479 dvdd.n478 0.429489
R3708 dvdd.n258 dvdd.n116 0.42139
R3709 dvdd.n356 dvdd.n300 0.410826
R3710 dvdd.n349 dvdd.n302 0.410826
R3711 dvdd.n393 dvdd.n320 0.410826
R3712 dvdd.n382 dvdd.n381 0.410826
R3713 dvdd.n454 dvdd.n453 0.383652
R3714 dvdd.n460 dvdd.n454 0.383652
R3715 dvdd.n430 dvdd.n428 0.383652
R3716 dvdd.n483 dvdd.n428 0.383652
R3717 dvdd.n437 dvdd.n432 0.383652
R3718 dvdd.n438 dvdd.n437 0.383652
R3719 dvdd.n475 dvdd.n433 0.383652
R3720 dvdd.n472 dvdd.n433 0.383652
R3721 dvdd.n435 dvdd.n434 0.383652
R3722 dvdd.n443 dvdd.n435 0.383652
R3723 dvdd.n471 dvdd.n444 0.383652
R3724 dvdd.n468 dvdd.n444 0.383652
R3725 dvdd.n446 dvdd.n445 0.383652
R3726 dvdd.n447 dvdd.n446 0.383652
R3727 dvdd.n467 dvdd.n448 0.383652
R3728 dvdd.n464 dvdd.n448 0.383652
R3729 dvdd.n450 dvdd.n449 0.383652
R3730 dvdd.n451 dvdd.n450 0.383652
R3731 dvdd.n463 dvdd.n452 0.383652
R3732 dvdd.n279 dvdd.n278 0.383652
R3733 dvdd.n278 dvdd.n277 0.383652
R3734 dvdd.n511 dvdd.n510 0.383652
R3735 dvdd.n510 dvdd.n509 0.383652
R3736 dvdd.n313 dvdd.n312 0.383652
R3737 dvdd.n314 dvdd.n313 0.383652
R3738 dvdd.n330 dvdd.n329 0.383652
R3739 dvdd.n377 dvdd.n324 0.383652
R3740 dvdd.n327 dvdd.n324 0.383652
R3741 dvdd.n378 dvdd.n323 0.383652
R3742 dvdd.n323 dvdd.n322 0.383652
R3743 dvdd.n373 dvdd.n326 0.383652
R3744 dvdd.n376 dvdd.n326 0.383652
R3745 dvdd.n333 dvdd.n332 0.383652
R3746 dvdd.n332 dvdd.n331 0.383652
R3747 dvdd.n369 dvdd.n334 0.383652
R3748 dvdd.n372 dvdd.n334 0.383652
R3749 dvdd.n337 dvdd.n336 0.383652
R3750 dvdd.n336 dvdd.n335 0.383652
R3751 dvdd.n365 dvdd.n338 0.383652
R3752 dvdd.n368 dvdd.n338 0.383652
R3753 dvdd.n341 dvdd.n340 0.383652
R3754 dvdd.n340 dvdd.n339 0.383652
R3755 dvdd.n361 dvdd.n342 0.383652
R3756 dvdd.n364 dvdd.n342 0.383652
R3757 dvdd.n345 dvdd.n344 0.383652
R3758 dvdd.n344 dvdd.n343 0.383652
R3759 dvdd.n353 dvdd.n346 0.383652
R3760 dvdd.n360 dvdd.n346 0.383652
R3761 dvdd.n354 dvdd.n348 0.383652
R3762 dvdd.n359 dvdd.n348 0.383652
R3763 dvdd.n351 dvdd.n350 0.383652
R3764 dvdd.n416 dvdd.n299 0.383652
R3765 dvdd.n413 dvdd.n299 0.383652
R3766 dvdd.n301 dvdd.n300 0.383652
R3767 dvdd.n302 dvdd.n301 0.383652
R3768 dvdd.n412 dvdd.n303 0.383652
R3769 dvdd.n409 dvdd.n303 0.383652
R3770 dvdd.n305 dvdd.n304 0.383652
R3771 dvdd.n306 dvdd.n305 0.383652
R3772 dvdd.n408 dvdd.n307 0.383652
R3773 dvdd.n405 dvdd.n307 0.383652
R3774 dvdd.n309 dvdd.n308 0.383652
R3775 dvdd.n310 dvdd.n309 0.383652
R3776 dvdd.n404 dvdd.n311 0.383652
R3777 dvdd.n400 dvdd.n311 0.383652
R3778 dvdd.n318 dvdd.n317 0.383652
R3779 dvdd.n394 dvdd.n318 0.383652
R3780 dvdd.n400 dvdd.n397 0.383652
R3781 dvdd.n397 dvdd.n396 0.383652
R3782 dvdd.n393 dvdd.n319 0.383652
R3783 dvdd.n382 dvdd.n319 0.383652
R3784 dvdd.n383 dvdd.n316 0.383652
R3785 dvdd.n390 dvdd.n383 0.383652
R3786 dvdd.n385 dvdd.n384 0.383652
R3787 dvdd.n389 dvdd.n385 0.383652
R3788 dvdd.n501 dvdd.n284 0.383652
R3789 dvdd.n387 dvdd.n284 0.383652
R3790 dvdd.n502 dvdd.n283 0.383652
R3791 dvdd.n283 dvdd.n282 0.383652
R3792 dvdd.n497 dvdd.n286 0.383652
R3793 dvdd.n500 dvdd.n286 0.383652
R3794 dvdd.n492 dvdd.n291 0.383652
R3795 dvdd.n399 dvdd.n291 0.383652
R3796 dvdd.n399 dvdd.n398 0.383652
R3797 dvdd.n398 dvdd.n287 0.383652
R3798 dvdd.n495 dvdd.n494 0.383652
R3799 dvdd.n496 dvdd.n495 0.383652
R3800 dvdd.n293 dvdd.n292 0.383652
R3801 dvdd.n491 dvdd.n292 0.383652
R3802 dvdd.n487 dvdd.n295 0.383652
R3803 dvdd.n297 dvdd.n295 0.383652
R3804 dvdd.n488 dvdd.n294 0.383652
R3805 dvdd.n294 dvdd.n290 0.383652
R3806 dvdd.n420 dvdd.n416 0.373755
R3807 dvdd.n484 dvdd.n427 0.373227
R3808 dvdd.n400 dvdd.n399 0.373
R3809 dvdd.n461 dvdd.n460 0.351043
R3810 dvdd.n474 dvdd.n434 0.351043
R3811 dvdd.n475 dvdd.n474 0.351043
R3812 dvdd.n473 dvdd.n443 0.351043
R3813 dvdd.n473 dvdd.n472 0.351043
R3814 dvdd.n470 dvdd.n445 0.351043
R3815 dvdd.n471 dvdd.n470 0.351043
R3816 dvdd.n469 dvdd.n447 0.351043
R3817 dvdd.n469 dvdd.n468 0.351043
R3818 dvdd.n466 dvdd.n449 0.351043
R3819 dvdd.n467 dvdd.n466 0.351043
R3820 dvdd.n465 dvdd.n451 0.351043
R3821 dvdd.n465 dvdd.n464 0.351043
R3822 dvdd.n462 dvdd.n453 0.351043
R3823 dvdd.n463 dvdd.n462 0.351043
R3824 dvdd.n328 dvdd.n327 0.351043
R3825 dvdd.n330 dvdd.n325 0.351043
R3826 dvdd.n377 dvdd.n325 0.351043
R3827 dvdd.n375 dvdd.n331 0.351043
R3828 dvdd.n376 dvdd.n375 0.351043
R3829 dvdd.n374 dvdd.n333 0.351043
R3830 dvdd.n374 dvdd.n373 0.351043
R3831 dvdd.n371 dvdd.n335 0.351043
R3832 dvdd.n372 dvdd.n371 0.351043
R3833 dvdd.n370 dvdd.n337 0.351043
R3834 dvdd.n370 dvdd.n369 0.351043
R3835 dvdd.n367 dvdd.n339 0.351043
R3836 dvdd.n368 dvdd.n367 0.351043
R3837 dvdd.n366 dvdd.n341 0.351043
R3838 dvdd.n366 dvdd.n365 0.351043
R3839 dvdd.n363 dvdd.n343 0.351043
R3840 dvdd.n364 dvdd.n363 0.351043
R3841 dvdd.n362 dvdd.n345 0.351043
R3842 dvdd.n362 dvdd.n361 0.351043
R3843 dvdd.n350 dvdd.n347 0.351043
R3844 dvdd.n360 dvdd.n347 0.351043
R3845 dvdd.n353 dvdd.n352 0.351043
R3846 dvdd.n415 dvdd.n300 0.351043
R3847 dvdd.n416 dvdd.n415 0.351043
R3848 dvdd.n414 dvdd.n302 0.351043
R3849 dvdd.n414 dvdd.n413 0.351043
R3850 dvdd.n411 dvdd.n304 0.351043
R3851 dvdd.n412 dvdd.n411 0.351043
R3852 dvdd.n410 dvdd.n306 0.351043
R3853 dvdd.n410 dvdd.n409 0.351043
R3854 dvdd.n407 dvdd.n308 0.351043
R3855 dvdd.n408 dvdd.n407 0.351043
R3856 dvdd.n406 dvdd.n310 0.351043
R3857 dvdd.n406 dvdd.n405 0.351043
R3858 dvdd.n403 dvdd.n312 0.351043
R3859 dvdd.n404 dvdd.n403 0.351043
R3860 dvdd.n402 dvdd.n314 0.351043
R3861 dvdd.n317 dvdd.n315 0.351043
R3862 dvdd.n395 dvdd.n394 0.351043
R3863 dvdd.n396 dvdd.n395 0.351043
R3864 dvdd.n393 dvdd.n392 0.351043
R3865 dvdd.n392 dvdd.n316 0.351043
R3866 dvdd.n391 dvdd.n382 0.351043
R3867 dvdd.n391 dvdd.n390 0.351043
R3868 dvdd.n389 dvdd.n388 0.351043
R3869 dvdd.n388 dvdd.n387 0.351043
R3870 dvdd.n384 dvdd.n285 0.351043
R3871 dvdd.n501 dvdd.n285 0.351043
R3872 dvdd.n498 dvdd.n497 0.351043
R3873 dvdd.n499 dvdd.n287 0.351043
R3874 dvdd.n500 dvdd.n499 0.351043
R3875 dvdd.n496 dvdd.n289 0.351043
R3876 dvdd.n493 dvdd.n492 0.351043
R3877 dvdd.n494 dvdd.n493 0.351043
R3878 dvdd.n491 dvdd.n490 0.351043
R3879 dvdd.n490 dvdd.n290 0.351043
R3880 dvdd.n489 dvdd.n293 0.351043
R3881 dvdd.n489 dvdd.n488 0.351043
R3882 dvdd.n507 dvdd.n506 0.307565
R3883 dvdd.n402 dvdd.n401 0.288543
R3884 dvdd.n401 dvdd.n315 0.288543
R3885 dvdd.n498 dvdd.n288 0.288543
R3886 dvdd.n289 dvdd.n288 0.288543
R3887 dvdd.n439 dvdd.n436 0.263321
R3888 dvdd.n442 dvdd.n436 0.263321
R3889 dvdd.n431 dvdd.n429 0.263321
R3890 dvdd.n456 dvdd.n455 0.263321
R3891 dvdd.n459 dvdd.n455 0.263321
R3892 dvdd.n514 dvdd.n513 0.263321
R3893 dvdd.n515 dvdd.n514 0.263321
R3894 dvdd.n281 dvdd.n280 0.263321
R3895 dvdd.n506 dvdd.n281 0.263321
R3896 dvdd.n480 dvdd.n431 0.226462
R3897 dvdd.n356 dvdd.n355 0.2055
R3898 dvdd.n355 dvdd.n349 0.2055
R3899 dvdd.n321 dvdd.n320 0.20347
R3900 dvdd.n381 dvdd.n321 0.20347
R3901 dvdd.n252 dvdd.n103 0.198679
R3902 dvdd.n663 dvdd 0.177824
R3903 dvdd.n663 dvdd.n49 0.170597
R3904 dvdd.n509 dvdd.n507 0.163543
R3905 dvdd.n665 dvdd 0.155803
R3906 dvdd.n666 dvdd 0.155803
R3907 dvdd.n667 dvdd 0.155803
R3908 dvdd.n387 dvdd.n386 0.141804
R3909 dvdd.n484 dvdd.n298 0.1255
R3910 dvdd.n479 dvdd.n432 0.0646892
R3911 dvdd.n478 dvdd.n476 0.0616026
R3912 dvdd.n421 dvdd.n420 0.0612215
R3913 dvdd.n430 dvdd.n50 0.0579324
R3914 dvdd.n480 dvdd.n479 0.0556802
R3915 dvdd.n427 dvdd.n50 0.0556802
R3916 dvdd.n46 dvdd.n45 0.0556724
R3917 dvdd.n34 dvdd.n33 0.0556724
R3918 dvdd.n22 dvdd.n21 0.0556724
R3919 dvdd.n10 dvdd.n9 0.0556724
R3920 dvdd.n662 dvdd.n50 0.0414555
R3921 dvdd dvdd.n47 0.0390101
R3922 dvdd dvdd.n35 0.0390101
R3923 dvdd dvdd.n23 0.0390101
R3924 dvdd dvdd.n11 0.0390101
R3925 dvdd.n269 dvdd.n260 0.0329873
R3926 dvdd.n662 dvdd.n661 0.0196358
R3927 dvdd.n476 dvdd 0.0171413
R3928 dvdd.n663 dvdd.n662 0.0165004
R3929 dvdd.n427 dvdd.n426 0.0162658
R3930 dvdd.n479 dvdd.n49 0.0139654
R3931 dvdd.n401 dvdd.n400 0.012
R3932 dvdd.n399 dvdd.n288 0.012
R3933 dvdd.n664 dvdd 0.0109536
R3934 dvdd.n423 dvdd.n50 0.00386852
R3935 dvdd.n425 dvdd.n424 0.00189736
R3936 dvdd.n424 dvdd.n423 0.000668426
R3937 comp_hyst_0.net3.t8 comp_hyst_0.net3.n1 242.409
R3938 comp_hyst_0.net3.n21 comp_hyst_0.net3.n1 1.7055
R3939 comp_hyst_0.net3.n1 comp_hyst_0.net3.n0 6.59063
R3940 comp_hyst_0.net3.n19 comp_hyst_0.net3.n20 0.244833
R3941 comp_hyst_0.net3.n21 comp_hyst_0.net3.n19 0.190675
R3942 comp_hyst_0.net3.n18 comp_hyst_0.net3.n21 0.194873
R3943 comp_hyst_0.net3.n10 comp_hyst_0.net3.n18 0.0950311
R3944 comp_hyst_0.net3.n9 comp_hyst_0.net3.n10 0.0472345
R3945 comp_hyst_0.net3 comp_hyst_0.net3.n9 0.087065
R3946 comp_hyst_0.net3.n20 comp_hyst_0.net3.t0 85.4116
R3947 comp_hyst_0.net3.n20 comp_hyst_0.net3.t1 85.24
R3948 comp_hyst_0.net3.n19 comp_hyst_0.net3.t12 86.0843
R3949 comp_hyst_0.net3.n12 comp_hyst_0.net3.n11 0.0905
R3950 comp_hyst_0.net3.n17 comp_hyst_0.net3.n12 5.44738
R3951 comp_hyst_0.net3.n18 comp_hyst_0.net3.n17 5.41956
R3952 comp_hyst_0.net3.n17 comp_hyst_0.net3.t13 6.00662
R3953 comp_hyst_0.net3.n16 comp_hyst_0.net3.t13 6.00662
R3954 comp_hyst_0.net3.n15 comp_hyst_0.net3.n13 0.0905
R3955 comp_hyst_0.net3.n16 comp_hyst_0.net3.n15 5.44738
R3956 comp_hyst_0.net3.n10 comp_hyst_0.net3.n16 5.41956
R3957 comp_hyst_0.net3.n15 comp_hyst_0.net3.t11 11.4535
R3958 comp_hyst_0.net3.n12 comp_hyst_0.net3.t11 11.4535
R3959 comp_hyst_0.net3.n13 comp_hyst_0.net3.n14 3.61579
R3960 comp_hyst_0.net3.n11 comp_hyst_0.net3.n14 3.61579
R3961 comp_hyst_0.net3.n11 comp_hyst_0.net3.t4 5.91616
R3962 comp_hyst_0.net3.n13 comp_hyst_0.net3.t4 5.91616
R3963 comp_hyst_0.net3.n14 comp_hyst_0.net3.t5 228.215
R3964 comp_hyst_0.net3.n3 comp_hyst_0.net3.n2 0.0905
R3965 comp_hyst_0.net3.n8 comp_hyst_0.net3.n3 5.44738
R3966 comp_hyst_0.net3.n9 comp_hyst_0.net3.n8 5.41956
R3967 comp_hyst_0.net3.n8 comp_hyst_0.net3.t10 6.00662
R3968 comp_hyst_0.net3.n7 comp_hyst_0.net3.t10 6.00662
R3969 comp_hyst_0.net3.n6 comp_hyst_0.net3.n4 0.0905
R3970 comp_hyst_0.net3.n7 comp_hyst_0.net3.n6 5.44738
R3971 comp_hyst_0.net3 comp_hyst_0.net3.n7 5.42753
R3972 comp_hyst_0.net3.n6 comp_hyst_0.net3.t9 11.4535
R3973 comp_hyst_0.net3.n3 comp_hyst_0.net3.t9 11.4535
R3974 comp_hyst_0.net3.n4 comp_hyst_0.net3.n5 3.61579
R3975 comp_hyst_0.net3.n2 comp_hyst_0.net3.n5 3.61579
R3976 comp_hyst_0.net3.n2 comp_hyst_0.net3.t6 5.91616
R3977 comp_hyst_0.net3.n4 comp_hyst_0.net3.t6 5.91616
R3978 comp_hyst_0.net3.n5 comp_hyst_0.net3.t7 228.215
R3979 comp_hyst_0.net3.n0 comp_hyst_0.net3.t3 231.423
R3980 comp_hyst_0.net3.n0 comp_hyst_0.net3.t2 232.41
R3981 level_shifter_3.in_b.n0 level_shifter_3.in_b.t1 83.7172
R3982 level_shifter_3.in_b.n0 level_shifter_3.in_b.t0 229.644
R3983 level_shifter_3.in_b level_shifter_3.in_b.n0 5.2032
R3984 level_shifter_3.in_b level_shifter_3.in_b.t2 21.9226
R3985 multiplexer_0.vtrip_3.n0 multiplexer_0.vtrip_3.t1 41.2565
R3986 multiplexer_0.vtrip_3.n1 multiplexer_0.vtrip_3.n0 5.29988
R3987 multiplexer_0.vtrip_3.n1 multiplexer_0.vtrip_3.t2 16.8956
R3988 multiplexer_0.vtrip_3 multiplexer_0.vtrip_3.n1 1.62926
R3989 multiplexer_0.vtrip_3 multiplexer_0.vtrip_3.n2 0.171398
R3990 multiplexer_0.vtrip_3.n2 multiplexer_0.vtrip_3.n3 1.3589
R3991 multiplexer_0.vtrip_3.t4 multiplexer_0.vtrip_3.n3 97.296
R3992 multiplexer_0.vtrip_3.n3 multiplexer_0.vtrip_3 4.98306
R3993 multiplexer_0.vtrip_3.t5 multiplexer_0.vtrip_3 18.5516
R3994 multiplexer_0.vtrip_3.n2 multiplexer_0.vtrip_3 3.32193
R3995 multiplexer_0.vtrip_3 multiplexer_0.vtrip_3.t3 18.1873
R3996 multiplexer_0.vtrip_3.n0 multiplexer_0.vtrip_3.t0 227.385
R3997 a_n8362_4845.t0 a_n8362_4845.t1 21.2567
R3998 multiplexer_0.in_0110.n0 multiplexer_0.in_0110.t3 228.216
R3999 multiplexer_0.in_0110.n0 multiplexer_0.in_0110.t2 83.695
R4000 multiplexer_0.in_0110.n4 multiplexer_0.in_0110.t0 10.5295
R4001 multiplexer_0.in_0110.n4 multiplexer_0.in_0110.t1 10.5285
R4002 multiplexer_0.in_0110 multiplexer_0.in_0110.n3 4.51461
R4003 multiplexer_0.in_0110.n2 multiplexer_0.in_0110.n1 4.34635
R4004 multiplexer_0.in_0110.n1 multiplexer_0.in_0110.n0 1.5005
R4005 multiplexer_0.in_0110 multiplexer_0.in_0110.n4 0.872792
R4006 multiplexer_0.in_0110.n3 multiplexer_0.in_0110 0.177654
R4007 multiplexer_0.in_0110.n1 multiplexer_0.in_0110 0.104667
R4008 multiplexer_0.in_0110.n2 multiplexer_0.in_0110 0.0064902
R4009 multiplexer_0.in_0110.n3 multiplexer_0.in_0110.n2 0.00411538
R4010 a_n15874_8625.t0 a_n15874_8625.t1 21.2567
R4011 a_n12654_9003.t0 a_n12654_9003.t1 21.167
R4012 multiplexer_0.vtrip_2.n0 multiplexer_0.vtrip_2.t1 41.2565
R4013 multiplexer_0.vtrip_2.n1 multiplexer_0.vtrip_2.n0 5.29988
R4014 multiplexer_0.vtrip_2.n1 multiplexer_0.vtrip_2.t6 16.8956
R4015 multiplexer_0.vtrip_2 multiplexer_0.vtrip_2.n1 1.62926
R4016 multiplexer_0.vtrip_2 multiplexer_0.vtrip_2.n6 13.7934
R4017 multiplexer_0.vtrip_2 multiplexer_0.vtrip_2.n6 5.50552
R4018 multiplexer_0.vtrip_2.n6 multiplexer_0.vtrip_2.n5 2.31984
R4019 multiplexer_0.vtrip_2.n5 multiplexer_0.vtrip_2.t2 97.296
R4020 multiplexer_0.vtrip_2.n5 multiplexer_0.vtrip_2.n3 0.0893672
R4021 multiplexer_0.vtrip_2.n3 multiplexer_0.vtrip_2.n2 4.7173
R4022 multiplexer_0.vtrip_2.n2 multiplexer_0.vtrip_2 0.103039
R4023 multiplexer_0.vtrip_2.n3 multiplexer_0.vtrip_2 3.32193
R4024 multiplexer_0.vtrip_2 multiplexer_0.vtrip_2.n4 1.67907
R4025 multiplexer_0.vtrip_2.t3 multiplexer_0.vtrip_2.n4 16.8731
R4026 multiplexer_0.vtrip_2.n4 multiplexer_0.vtrip_2.t5 16.5088
R4027 multiplexer_0.vtrip_2.n2 multiplexer_0.vtrip_2 3.32193
R4028 multiplexer_0.vtrip_2.t4 multiplexer_0.vtrip_2 18.5516
R4029 multiplexer_0.vtrip_2 multiplexer_0.vtrip_2.t7 18.1873
R4030 multiplexer_0.vtrip_2.n0 multiplexer_0.vtrip_2.t0 227.385
R4031 a_n12118_9759.t0 a_n12118_9759.t1 21.2567
R4032 a_n8898_9381.t0 a_n8898_9381.t1 21.167
R4033 multiplexer_0.in_1100.n0 multiplexer_0.in_1100.t3 228.216
R4034 multiplexer_0.in_1100.n0 multiplexer_0.in_1100.t2 83.695
R4035 multiplexer_0.in_1100.n3 multiplexer_0.in_1100.t1 10.5739
R4036 multiplexer_0.in_1100.n3 multiplexer_0.in_1100.t0 10.5739
R4037 multiplexer_0.in_1100 multiplexer_0.in_1100.n3 2.20538
R4038 multiplexer_0.in_1100 multiplexer_0.in_1100.n0 1.60467
R4039 multiplexer_0.in_1100 multiplexer_0.in_1100.n2 0.9755
R4040 multiplexer_0.in_1100.n2 multiplexer_0.in_1100 0.471654
R4041 multiplexer_0.in_1100.n1 multiplexer_0.in_1100 0.414042
R4042 multiplexer_0.in_1100.n1 multiplexer_0.in_1100 0.0140417
R4043 multiplexer_0.in_1100.n2 multiplexer_0.in_1100.n1 0.0101154
R4044 multiplexer_0.in_1101.n0 multiplexer_0.in_1101.t0 228.216
R4045 multiplexer_0.in_1101.n0 multiplexer_0.in_1101.t1 83.695
R4046 multiplexer_0.in_1101.n3 multiplexer_0.in_1101.t2 10.5295
R4047 multiplexer_0.in_1101.n3 multiplexer_0.in_1101.t3 10.5285
R4048 multiplexer_0.in_1101 multiplexer_0.in_1101.n2 3.98817
R4049 multiplexer_0.in_1101 multiplexer_0.in_1101.n0 1.60467
R4050 multiplexer_0.in_1101 multiplexer_0.in_1101.n3 0.872792
R4051 multiplexer_0.in_1101.n2 multiplexer_0.in_1101 0.471654
R4052 multiplexer_0.in_1101.n1 multiplexer_0.in_1101 0.414042
R4053 multiplexer_0.in_1101.n1 multiplexer_0.in_1101 0.0140417
R4054 multiplexer_0.in_1101.n2 multiplexer_0.in_1101.n1 0.0101154
R4055 a_n15874_6357.t0 a_n15874_6357.t1 21.2567
R4056 a_n12654_5979.t0 a_n12654_5979.t1 21.167
R4057 vtrip[0].n2 vtrip[0].t2 99.4021
R4058 vtrip[0].n0 vtrip[0].t1 23.1698
R4059 vtrip[0].n1 vtrip[0].t3 17.7681
R4060 vtrip[0].n0 vtrip[0].t0 17.7475
R4061 vtrip[0].n2 vtrip[0] 5.62823
R4062 vtrip[0].n3 vtrip[0].n2 1.7055
R4063 vtrip[0].n1 vtrip[0].n0 0.572059
R4064 vtrip[0].n3 vtrip[0].n1 0.1139
R4065 vtrip[0] vtrip[0].n3 0.0378665
R4066 level_shifter_0.in_b.n0 level_shifter_0.in_b.t1 83.7172
R4067 level_shifter_0.in_b.n0 level_shifter_0.in_b.t0 229.644
R4068 level_shifter_0.in_b level_shifter_0.in_b.n0 5.2032
R4069 level_shifter_0.in_b level_shifter_0.in_b.t2 21.9226
R4070 multiplexer_0.trans_gate_m_32.in.t1 multiplexer_0.trans_gate_m_32.in.n0 228.216
R4071 multiplexer_0.trans_gate_m_32.in.n5 multiplexer_0.trans_gate_m_32.in.n0 1.5005
R4072 multiplexer_0.trans_gate_m_32.in.n0 multiplexer_0.trans_gate_m_32.in.t5 83.695
R4073 multiplexer_0.trans_gate_m_32.in multiplexer_0.trans_gate_m_32.in.n5 0.104667
R4074 multiplexer_0.trans_gate_m_32.in.n4 multiplexer_0.trans_gate_m_32.in.n5 0.459875
R4075 multiplexer_0.trans_gate_m_32.in multiplexer_0.trans_gate_m_32.in.n4 0.553625
R4076 multiplexer_0.trans_gate_m_32.in multiplexer_0.trans_gate_m_32.in.n1 1.60467
R4077 multiplexer_0.trans_gate_m_32.in.n4 multiplexer_0.trans_gate_m_32.in.n3 4.43682
R4078 multiplexer_0.trans_gate_m_32.in.n3 multiplexer_0.trans_gate_m_32.in.n2 1.5005
R4079 multiplexer_0.trans_gate_m_32.in multiplexer_0.trans_gate_m_32.in.n3 0.104667
R4080 multiplexer_0.trans_gate_m_32.in.n2 multiplexer_0.trans_gate_m_32.in.t2 83.695
R4081 multiplexer_0.trans_gate_m_32.in.n2 multiplexer_0.trans_gate_m_32.in.t4 228.216
R4082 multiplexer_0.trans_gate_m_32.in.n1 multiplexer_0.trans_gate_m_32.in.t0 83.695
R4083 multiplexer_0.trans_gate_m_32.in.n1 multiplexer_0.trans_gate_m_32.in.t3 228.216
R4084 multiplexer_0.trans_gate_m_37.out.t1 multiplexer_0.trans_gate_m_37.out.n0 228.216
R4085 multiplexer_0.trans_gate_m_37.out.n5 multiplexer_0.trans_gate_m_37.out.n0 1.5005
R4086 multiplexer_0.trans_gate_m_37.out.n0 multiplexer_0.trans_gate_m_37.out.t4 83.695
R4087 multiplexer_0.trans_gate_m_37.out multiplexer_0.trans_gate_m_37.out.n5 0.104667
R4088 multiplexer_0.trans_gate_m_37.out.n5 multiplexer_0.trans_gate_m_37.out.n4 5.41376
R4089 multiplexer_0.trans_gate_m_37.out.n2 multiplexer_0.trans_gate_m_37.out.n1 1.5005
R4090 multiplexer_0.trans_gate_m_37.out multiplexer_0.trans_gate_m_37.out.n2 0.104667
R4091 multiplexer_0.trans_gate_m_37.out.n4 multiplexer_0.trans_gate_m_37.out.n2 0.459875
R4092 multiplexer_0.trans_gate_m_37.out.n4 multiplexer_0.trans_gate_m_37.out 0.563
R4093 multiplexer_0.trans_gate_m_37.out multiplexer_0.trans_gate_m_37.out.n3 1.60467
R4094 multiplexer_0.trans_gate_m_37.out.n3 multiplexer_0.trans_gate_m_37.out.t3 83.695
R4095 multiplexer_0.trans_gate_m_37.out.n3 multiplexer_0.trans_gate_m_37.out.t2 228.216
R4096 multiplexer_0.trans_gate_m_37.out.n1 multiplexer_0.trans_gate_m_37.out.t0 83.695
R4097 multiplexer_0.trans_gate_m_37.out.n1 multiplexer_0.trans_gate_m_37.out.t5 228.216
R4098 avdd.n84 avdd.n78 1446.62
R4099 avdd.n81 avdd.n80 1446.62
R4100 avdd.n73 avdd.n67 1446.62
R4101 avdd.n70 avdd.n69 1446.62
R4102 avdd.n62 avdd.n56 1446.62
R4103 avdd.n59 avdd.n58 1446.62
R4104 avdd.n51 avdd.n45 1446.62
R4105 avdd.n48 avdd.n47 1446.62
R4106 avdd.n40 avdd.n34 1446.62
R4107 avdd.n37 avdd.n36 1446.62
R4108 avdd.n29 avdd.n23 1446.62
R4109 avdd.n26 avdd.n25 1446.62
R4110 avdd.n18 avdd.n12 1446.62
R4111 avdd.n15 avdd.n14 1446.62
R4112 avdd.n7 avdd.n1 1446.62
R4113 avdd.n4 avdd.n3 1446.62
R4114 avdd.n172 avdd.n166 1446.62
R4115 avdd.n169 avdd.n168 1446.62
R4116 avdd.n161 avdd.n155 1446.62
R4117 avdd.n158 avdd.n157 1446.62
R4118 avdd.n150 avdd.n144 1446.62
R4119 avdd.n147 avdd.n146 1446.62
R4120 avdd.n139 avdd.n133 1446.62
R4121 avdd.n136 avdd.n135 1446.62
R4122 avdd.n128 avdd.n122 1446.62
R4123 avdd.n125 avdd.n124 1446.62
R4124 avdd.n117 avdd.n111 1446.62
R4125 avdd.n114 avdd.n113 1446.62
R4126 avdd.n106 avdd.n100 1446.62
R4127 avdd.n103 avdd.n102 1446.62
R4128 avdd.n95 avdd.n89 1446.62
R4129 avdd.n92 avdd.n91 1446.62
R4130 avdd.n260 avdd.n254 1446.62
R4131 avdd.n257 avdd.n256 1446.62
R4132 avdd.n249 avdd.n243 1446.62
R4133 avdd.n246 avdd.n245 1446.62
R4134 avdd.n238 avdd.n232 1446.62
R4135 avdd.n235 avdd.n234 1446.62
R4136 avdd.n227 avdd.n221 1446.62
R4137 avdd.n224 avdd.n223 1446.62
R4138 avdd.n216 avdd.n210 1446.62
R4139 avdd.n213 avdd.n212 1446.62
R4140 avdd.n205 avdd.n199 1446.62
R4141 avdd.n202 avdd.n201 1446.62
R4142 avdd.n194 avdd.n188 1446.62
R4143 avdd.n191 avdd.n190 1446.62
R4144 avdd.n183 avdd.n177 1446.62
R4145 avdd.n180 avdd.n179 1446.62
R4146 avdd.n304 avdd.n298 1446.62
R4147 avdd.n301 avdd.n300 1446.62
R4148 avdd.n293 avdd.n287 1446.62
R4149 avdd.n290 avdd.n289 1446.62
R4150 avdd.n282 avdd.n276 1446.62
R4151 avdd.n279 avdd.n278 1446.62
R4152 avdd.n271 avdd.n265 1446.62
R4153 avdd.n268 avdd.n267 1446.62
R4154 avdd.n326 avdd.n319 1446.62
R4155 avdd.n326 avdd.n317 1446.62
R4156 avdd.n327 avdd.n311 1446.62
R4157 avdd.n327 avdd.n312 1446.62
R4158 avdd.n349 avdd.n342 1446.62
R4159 avdd.n349 avdd.n340 1446.62
R4160 avdd.n350 avdd.n334 1446.62
R4161 avdd.n350 avdd.n335 1446.62
R4162 avdd.n373 avdd.n366 1446.62
R4163 avdd.n373 avdd.n364 1446.62
R4164 avdd.n374 avdd.n358 1446.62
R4165 avdd.n374 avdd.n359 1446.62
R4166 avdd.n397 avdd.n390 1446.62
R4167 avdd.n397 avdd.n388 1446.62
R4168 avdd.n398 avdd.n382 1446.62
R4169 avdd.n398 avdd.n383 1446.62
R4170 avdd.n316 avdd.n314 910.034
R4171 avdd.n318 avdd.n314 910.034
R4172 avdd.n339 avdd.n337 910.034
R4173 avdd.n341 avdd.n337 910.034
R4174 avdd.n363 avdd.n361 910.034
R4175 avdd.n365 avdd.n361 910.034
R4176 avdd.n387 avdd.n385 910.034
R4177 avdd.n389 avdd.n385 910.034
R4178 avdd.n319 avdd.n318 536.587
R4179 avdd.n316 avdd.n311 536.587
R4180 avdd.n317 avdd.n316 536.587
R4181 avdd.n318 avdd.n312 536.587
R4182 avdd.n342 avdd.n341 536.587
R4183 avdd.n339 avdd.n334 536.587
R4184 avdd.n340 avdd.n339 536.587
R4185 avdd.n341 avdd.n335 536.587
R4186 avdd.n366 avdd.n365 536.587
R4187 avdd.n363 avdd.n358 536.587
R4188 avdd.n364 avdd.n363 536.587
R4189 avdd.n365 avdd.n359 536.587
R4190 avdd.n390 avdd.n389 536.587
R4191 avdd.n387 avdd.n382 536.587
R4192 avdd.n388 avdd.n387 536.587
R4193 avdd.n389 avdd.n383 536.587
R4194 avdd.n82 avdd.n78 410.803
R4195 avdd.n83 avdd.n80 410.803
R4196 avdd.n71 avdd.n67 410.803
R4197 avdd.n72 avdd.n69 410.803
R4198 avdd.n60 avdd.n56 410.803
R4199 avdd.n61 avdd.n58 410.803
R4200 avdd.n49 avdd.n45 410.803
R4201 avdd.n50 avdd.n47 410.803
R4202 avdd.n38 avdd.n34 410.803
R4203 avdd.n39 avdd.n36 410.803
R4204 avdd.n27 avdd.n23 410.803
R4205 avdd.n28 avdd.n25 410.803
R4206 avdd.n16 avdd.n12 410.803
R4207 avdd.n17 avdd.n14 410.803
R4208 avdd.n5 avdd.n1 410.803
R4209 avdd.n6 avdd.n3 410.803
R4210 avdd.n170 avdd.n166 410.803
R4211 avdd.n171 avdd.n168 410.803
R4212 avdd.n159 avdd.n155 410.803
R4213 avdd.n160 avdd.n157 410.803
R4214 avdd.n148 avdd.n144 410.803
R4215 avdd.n149 avdd.n146 410.803
R4216 avdd.n137 avdd.n133 410.803
R4217 avdd.n138 avdd.n135 410.803
R4218 avdd.n126 avdd.n122 410.803
R4219 avdd.n127 avdd.n124 410.803
R4220 avdd.n115 avdd.n111 410.803
R4221 avdd.n116 avdd.n113 410.803
R4222 avdd.n104 avdd.n100 410.803
R4223 avdd.n105 avdd.n102 410.803
R4224 avdd.n93 avdd.n89 410.803
R4225 avdd.n94 avdd.n91 410.803
R4226 avdd.n258 avdd.n254 410.803
R4227 avdd.n259 avdd.n256 410.803
R4228 avdd.n247 avdd.n243 410.803
R4229 avdd.n248 avdd.n245 410.803
R4230 avdd.n236 avdd.n232 410.803
R4231 avdd.n237 avdd.n234 410.803
R4232 avdd.n225 avdd.n221 410.803
R4233 avdd.n226 avdd.n223 410.803
R4234 avdd.n214 avdd.n210 410.803
R4235 avdd.n215 avdd.n212 410.803
R4236 avdd.n203 avdd.n199 410.803
R4237 avdd.n204 avdd.n201 410.803
R4238 avdd.n192 avdd.n188 410.803
R4239 avdd.n193 avdd.n190 410.803
R4240 avdd.n181 avdd.n177 410.803
R4241 avdd.n182 avdd.n179 410.803
R4242 avdd.n302 avdd.n298 410.803
R4243 avdd.n303 avdd.n300 410.803
R4244 avdd.n291 avdd.n287 410.803
R4245 avdd.n292 avdd.n289 410.803
R4246 avdd.n280 avdd.n276 410.803
R4247 avdd.n281 avdd.n278 410.803
R4248 avdd.n269 avdd.n265 410.803
R4249 avdd.n270 avdd.n267 410.803
R4250 avdd.t24 avdd.n313 314.628
R4251 avdd.t24 avdd.n315 314.628
R4252 avdd.t1 avdd.n336 314.628
R4253 avdd.t1 avdd.n338 314.628
R4254 avdd.t18 avdd.n360 314.628
R4255 avdd.t18 avdd.n362 314.628
R4256 avdd.t13 avdd.n384 314.628
R4257 avdd.t13 avdd.n386 314.628
R4258 avdd.n85 avdd.n79 281.601
R4259 avdd.n74 avdd.n68 281.601
R4260 avdd.n63 avdd.n57 281.601
R4261 avdd.n52 avdd.n46 281.601
R4262 avdd.n41 avdd.n35 281.601
R4263 avdd.n30 avdd.n24 281.601
R4264 avdd.n19 avdd.n13 281.601
R4265 avdd.n8 avdd.n2 281.601
R4266 avdd.n173 avdd.n167 281.601
R4267 avdd.n162 avdd.n156 281.601
R4268 avdd.n151 avdd.n145 281.601
R4269 avdd.n140 avdd.n134 281.601
R4270 avdd.n129 avdd.n123 281.601
R4271 avdd.n118 avdd.n112 281.601
R4272 avdd.n107 avdd.n101 281.601
R4273 avdd.n96 avdd.n90 281.601
R4274 avdd.n261 avdd.n255 281.601
R4275 avdd.n250 avdd.n244 281.601
R4276 avdd.n239 avdd.n233 281.601
R4277 avdd.n228 avdd.n222 281.601
R4278 avdd.n217 avdd.n211 281.601
R4279 avdd.n206 avdd.n200 281.601
R4280 avdd.n195 avdd.n189 281.601
R4281 avdd.n184 avdd.n178 281.601
R4282 avdd.n305 avdd.n299 281.601
R4283 avdd.n294 avdd.n288 281.601
R4284 avdd.n283 avdd.n277 281.601
R4285 avdd.n272 avdd.n266 281.601
R4286 avdd.n308 avdd.t27 227.845
R4287 avdd.n331 avdd.t2 227.845
R4288 avdd.n355 avdd.t39 227.845
R4289 avdd.n379 avdd.t32 227.845
R4290 avdd.n308 avdd.t25 227.345
R4291 avdd.n331 avdd.t29 227.345
R4292 avdd.n355 avdd.t19 227.345
R4293 avdd.n379 avdd.t14 227.345
R4294 avdd.n79 avdd.n77 217.418
R4295 avdd.n68 avdd.n66 217.418
R4296 avdd.n57 avdd.n55 217.418
R4297 avdd.n46 avdd.n44 217.418
R4298 avdd.n35 avdd.n33 217.418
R4299 avdd.n24 avdd.n22 217.418
R4300 avdd.n13 avdd.n11 217.418
R4301 avdd.n2 avdd.n0 217.418
R4302 avdd.n167 avdd.n165 217.418
R4303 avdd.n156 avdd.n154 217.418
R4304 avdd.n145 avdd.n143 217.418
R4305 avdd.n134 avdd.n132 217.418
R4306 avdd.n123 avdd.n121 217.418
R4307 avdd.n112 avdd.n110 217.418
R4308 avdd.n101 avdd.n99 217.418
R4309 avdd.n90 avdd.n88 217.418
R4310 avdd.n255 avdd.n253 217.418
R4311 avdd.n244 avdd.n242 217.418
R4312 avdd.n233 avdd.n231 217.418
R4313 avdd.n222 avdd.n220 217.418
R4314 avdd.n211 avdd.n209 217.418
R4315 avdd.n200 avdd.n198 217.418
R4316 avdd.n189 avdd.n187 217.418
R4317 avdd.n178 avdd.n176 217.418
R4318 avdd.n299 avdd.n297 217.418
R4319 avdd.n288 avdd.n286 217.418
R4320 avdd.n277 avdd.n275 217.418
R4321 avdd.n266 avdd.n264 217.418
R4322 avdd.n86 avdd.n85 205.571
R4323 avdd.n75 avdd.n74 205.571
R4324 avdd.n64 avdd.n63 205.571
R4325 avdd.n53 avdd.n52 205.571
R4326 avdd.n42 avdd.n41 205.571
R4327 avdd.n31 avdd.n30 205.571
R4328 avdd.n20 avdd.n19 205.571
R4329 avdd.n9 avdd.n8 205.571
R4330 avdd.n174 avdd.n173 205.571
R4331 avdd.n163 avdd.n162 205.571
R4332 avdd.n152 avdd.n151 205.571
R4333 avdd.n141 avdd.n140 205.571
R4334 avdd.n130 avdd.n129 205.571
R4335 avdd.n119 avdd.n118 205.571
R4336 avdd.n108 avdd.n107 205.571
R4337 avdd.n97 avdd.n96 205.571
R4338 avdd.n262 avdd.n261 205.571
R4339 avdd.n251 avdd.n250 205.571
R4340 avdd.n240 avdd.n239 205.571
R4341 avdd.n229 avdd.n228 205.571
R4342 avdd.n218 avdd.n217 205.571
R4343 avdd.n207 avdd.n206 205.571
R4344 avdd.n196 avdd.n195 205.571
R4345 avdd.n185 avdd.n184 205.571
R4346 avdd.n306 avdd.n305 205.571
R4347 avdd.n295 avdd.n294 205.571
R4348 avdd.n284 avdd.n283 205.571
R4349 avdd.n273 avdd.n272 205.571
R4350 avdd.n322 avdd.n321 174.306
R4351 avdd.n323 avdd.n322 174.306
R4352 avdd.n345 avdd.n344 174.306
R4353 avdd.n346 avdd.n345 174.306
R4354 avdd.n369 avdd.n368 174.306
R4355 avdd.n370 avdd.n369 174.306
R4356 avdd.n393 avdd.n392 174.306
R4357 avdd.n394 avdd.n393 174.306
R4358 avdd.n328 avdd.n310 132.73
R4359 avdd.n351 avdd.n333 132.73
R4360 avdd.n375 avdd.n357 132.73
R4361 avdd.n399 avdd.n381 132.73
R4362 avdd.n329 avdd.n309 132.674
R4363 avdd.n352 avdd.n332 132.674
R4364 avdd.n376 avdd.n356 132.674
R4365 avdd.n400 avdd.n380 132.674
R4366 avdd.n86 avdd.n77 117.996
R4367 avdd.n75 avdd.n66 117.996
R4368 avdd.n64 avdd.n55 117.996
R4369 avdd.n53 avdd.n44 117.996
R4370 avdd.n42 avdd.n33 117.996
R4371 avdd.n31 avdd.n22 117.996
R4372 avdd.n20 avdd.n11 117.996
R4373 avdd.n9 avdd.n0 117.996
R4374 avdd.n174 avdd.n165 117.996
R4375 avdd.n163 avdd.n154 117.996
R4376 avdd.n152 avdd.n143 117.996
R4377 avdd.n141 avdd.n132 117.996
R4378 avdd.n130 avdd.n121 117.996
R4379 avdd.n119 avdd.n110 117.996
R4380 avdd.n108 avdd.n99 117.996
R4381 avdd.n97 avdd.n88 117.996
R4382 avdd.n262 avdd.n253 117.996
R4383 avdd.n251 avdd.n242 117.996
R4384 avdd.n240 avdd.n231 117.996
R4385 avdd.n229 avdd.n220 117.996
R4386 avdd.n218 avdd.n209 117.996
R4387 avdd.n207 avdd.n198 117.996
R4388 avdd.n196 avdd.n187 117.996
R4389 avdd.n185 avdd.n176 117.996
R4390 avdd.n306 avdd.n297 117.996
R4391 avdd.n295 avdd.n286 117.996
R4392 avdd.n284 avdd.n275 117.996
R4393 avdd.n273 avdd.n264 117.996
R4394 avdd.n325 avdd.n320 117.746
R4395 avdd.n325 avdd.n324 117.746
R4396 avdd.n348 avdd.n343 117.746
R4397 avdd.n348 avdd.n347 117.746
R4398 avdd.n372 avdd.n367 117.746
R4399 avdd.n372 avdd.n371 117.746
R4400 avdd.n396 avdd.n391 117.746
R4401 avdd.n396 avdd.n395 117.746
R4402 avdd.n321 avdd.n320 107.294
R4403 avdd.n323 avdd.n310 107.294
R4404 avdd.n324 avdd.n323 107.294
R4405 avdd.n321 avdd.n309 107.294
R4406 avdd.n344 avdd.n343 107.294
R4407 avdd.n346 avdd.n333 107.294
R4408 avdd.n347 avdd.n346 107.294
R4409 avdd.n344 avdd.n332 107.294
R4410 avdd.n368 avdd.n367 107.294
R4411 avdd.n370 avdd.n357 107.294
R4412 avdd.n371 avdd.n370 107.294
R4413 avdd.n368 avdd.n356 107.294
R4414 avdd.n392 avdd.n391 107.294
R4415 avdd.n394 avdd.n381 107.294
R4416 avdd.n395 avdd.n394 107.294
R4417 avdd.n392 avdd.n380 107.294
R4418 avdd.n80 avdd.n79 26.4291
R4419 avdd.n86 avdd.n78 26.4291
R4420 avdd.n69 avdd.n68 26.4291
R4421 avdd.n75 avdd.n67 26.4291
R4422 avdd.n58 avdd.n57 26.4291
R4423 avdd.n64 avdd.n56 26.4291
R4424 avdd.n47 avdd.n46 26.4291
R4425 avdd.n53 avdd.n45 26.4291
R4426 avdd.n36 avdd.n35 26.4291
R4427 avdd.n42 avdd.n34 26.4291
R4428 avdd.n25 avdd.n24 26.4291
R4429 avdd.n31 avdd.n23 26.4291
R4430 avdd.n14 avdd.n13 26.4291
R4431 avdd.n20 avdd.n12 26.4291
R4432 avdd.n3 avdd.n2 26.4291
R4433 avdd.n9 avdd.n1 26.4291
R4434 avdd.n168 avdd.n167 26.4291
R4435 avdd.n174 avdd.n166 26.4291
R4436 avdd.n157 avdd.n156 26.4291
R4437 avdd.n163 avdd.n155 26.4291
R4438 avdd.n146 avdd.n145 26.4291
R4439 avdd.n152 avdd.n144 26.4291
R4440 avdd.n135 avdd.n134 26.4291
R4441 avdd.n141 avdd.n133 26.4291
R4442 avdd.n124 avdd.n123 26.4291
R4443 avdd.n130 avdd.n122 26.4291
R4444 avdd.n113 avdd.n112 26.4291
R4445 avdd.n119 avdd.n111 26.4291
R4446 avdd.n102 avdd.n101 26.4291
R4447 avdd.n108 avdd.n100 26.4291
R4448 avdd.n91 avdd.n90 26.4291
R4449 avdd.n97 avdd.n89 26.4291
R4450 avdd.n256 avdd.n255 26.4291
R4451 avdd.n262 avdd.n254 26.4291
R4452 avdd.n245 avdd.n244 26.4291
R4453 avdd.n251 avdd.n243 26.4291
R4454 avdd.n234 avdd.n233 26.4291
R4455 avdd.n240 avdd.n232 26.4291
R4456 avdd.n223 avdd.n222 26.4291
R4457 avdd.n229 avdd.n221 26.4291
R4458 avdd.n212 avdd.n211 26.4291
R4459 avdd.n218 avdd.n210 26.4291
R4460 avdd.n201 avdd.n200 26.4291
R4461 avdd.n207 avdd.n199 26.4291
R4462 avdd.n190 avdd.n189 26.4291
R4463 avdd.n196 avdd.n188 26.4291
R4464 avdd.n179 avdd.n178 26.4291
R4465 avdd.n185 avdd.n177 26.4291
R4466 avdd.n300 avdd.n299 26.4291
R4467 avdd.n306 avdd.n298 26.4291
R4468 avdd.n289 avdd.n288 26.4291
R4469 avdd.n295 avdd.n287 26.4291
R4470 avdd.n278 avdd.n277 26.4291
R4471 avdd.n284 avdd.n276 26.4291
R4472 avdd.n267 avdd.n266 26.4291
R4473 avdd.n273 avdd.n265 26.4291
R4474 avdd.n320 avdd.n317 26.4291
R4475 avdd.n317 avdd.n313 26.4291
R4476 avdd.n312 avdd.n310 26.4291
R4477 avdd.n315 avdd.n312 26.4291
R4478 avdd.n324 avdd.n319 26.4291
R4479 avdd.n319 avdd.n315 26.4291
R4480 avdd.n311 avdd.n309 26.4291
R4481 avdd.n313 avdd.n311 26.4291
R4482 avdd.n343 avdd.n340 26.4291
R4483 avdd.n340 avdd.n336 26.4291
R4484 avdd.n335 avdd.n333 26.4291
R4485 avdd.n338 avdd.n335 26.4291
R4486 avdd.n347 avdd.n342 26.4291
R4487 avdd.n342 avdd.n338 26.4291
R4488 avdd.n334 avdd.n332 26.4291
R4489 avdd.n336 avdd.n334 26.4291
R4490 avdd.n367 avdd.n364 26.4291
R4491 avdd.n364 avdd.n360 26.4291
R4492 avdd.n359 avdd.n357 26.4291
R4493 avdd.n362 avdd.n359 26.4291
R4494 avdd.n371 avdd.n366 26.4291
R4495 avdd.n366 avdd.n362 26.4291
R4496 avdd.n358 avdd.n356 26.4291
R4497 avdd.n360 avdd.n358 26.4291
R4498 avdd.n391 avdd.n388 26.4291
R4499 avdd.n388 avdd.n384 26.4291
R4500 avdd.n383 avdd.n381 26.4291
R4501 avdd.n386 avdd.n383 26.4291
R4502 avdd.n395 avdd.n390 26.4291
R4503 avdd.n390 avdd.n386 26.4291
R4504 avdd.n382 avdd.n380 26.4291
R4505 avdd.n384 avdd.n382 26.4291
R4506 avdd.n81 avdd.n77 16.8187
R4507 avdd.n85 avdd.n84 16.8187
R4508 avdd.n70 avdd.n66 16.8187
R4509 avdd.n74 avdd.n73 16.8187
R4510 avdd.n59 avdd.n55 16.8187
R4511 avdd.n63 avdd.n62 16.8187
R4512 avdd.n48 avdd.n44 16.8187
R4513 avdd.n52 avdd.n51 16.8187
R4514 avdd.n37 avdd.n33 16.8187
R4515 avdd.n41 avdd.n40 16.8187
R4516 avdd.n26 avdd.n22 16.8187
R4517 avdd.n30 avdd.n29 16.8187
R4518 avdd.n15 avdd.n11 16.8187
R4519 avdd.n19 avdd.n18 16.8187
R4520 avdd.n4 avdd.n0 16.8187
R4521 avdd.n8 avdd.n7 16.8187
R4522 avdd.n169 avdd.n165 16.8187
R4523 avdd.n173 avdd.n172 16.8187
R4524 avdd.n158 avdd.n154 16.8187
R4525 avdd.n162 avdd.n161 16.8187
R4526 avdd.n147 avdd.n143 16.8187
R4527 avdd.n151 avdd.n150 16.8187
R4528 avdd.n136 avdd.n132 16.8187
R4529 avdd.n140 avdd.n139 16.8187
R4530 avdd.n125 avdd.n121 16.8187
R4531 avdd.n129 avdd.n128 16.8187
R4532 avdd.n114 avdd.n110 16.8187
R4533 avdd.n118 avdd.n117 16.8187
R4534 avdd.n103 avdd.n99 16.8187
R4535 avdd.n107 avdd.n106 16.8187
R4536 avdd.n92 avdd.n88 16.8187
R4537 avdd.n96 avdd.n95 16.8187
R4538 avdd.n257 avdd.n253 16.8187
R4539 avdd.n261 avdd.n260 16.8187
R4540 avdd.n246 avdd.n242 16.8187
R4541 avdd.n250 avdd.n249 16.8187
R4542 avdd.n235 avdd.n231 16.8187
R4543 avdd.n239 avdd.n238 16.8187
R4544 avdd.n224 avdd.n220 16.8187
R4545 avdd.n228 avdd.n227 16.8187
R4546 avdd.n213 avdd.n209 16.8187
R4547 avdd.n217 avdd.n216 16.8187
R4548 avdd.n202 avdd.n198 16.8187
R4549 avdd.n206 avdd.n205 16.8187
R4550 avdd.n191 avdd.n187 16.8187
R4551 avdd.n195 avdd.n194 16.8187
R4552 avdd.n180 avdd.n176 16.8187
R4553 avdd.n184 avdd.n183 16.8187
R4554 avdd.n301 avdd.n297 16.8187
R4555 avdd.n305 avdd.n304 16.8187
R4556 avdd.n290 avdd.n286 16.8187
R4557 avdd.n294 avdd.n293 16.8187
R4558 avdd.n279 avdd.n275 16.8187
R4559 avdd.n283 avdd.n282 16.8187
R4560 avdd.n268 avdd.n264 16.8187
R4561 avdd.n272 avdd.n271 16.8187
R4562 avdd.n326 avdd.n325 16.8187
R4563 avdd.t24 avdd.n326 16.8187
R4564 avdd.n322 avdd.n314 16.8187
R4565 avdd.t24 avdd.n314 16.8187
R4566 avdd.n328 avdd.n327 16.8187
R4567 avdd.n327 avdd.t24 16.8187
R4568 avdd.n349 avdd.n348 16.8187
R4569 avdd.t1 avdd.n349 16.8187
R4570 avdd.n345 avdd.n337 16.8187
R4571 avdd.t1 avdd.n337 16.8187
R4572 avdd.n351 avdd.n350 16.8187
R4573 avdd.n350 avdd.t1 16.8187
R4574 avdd.n373 avdd.n372 16.8187
R4575 avdd.t18 avdd.n373 16.8187
R4576 avdd.n369 avdd.n361 16.8187
R4577 avdd.t18 avdd.n361 16.8187
R4578 avdd.n375 avdd.n374 16.8187
R4579 avdd.n374 avdd.t18 16.8187
R4580 avdd.n397 avdd.n396 16.8187
R4581 avdd.t13 avdd.n397 16.8187
R4582 avdd.n393 avdd.n385 16.8187
R4583 avdd.t13 avdd.n385 16.8187
R4584 avdd.n399 avdd.n398 16.8187
R4585 avdd.n398 avdd.t13 16.8187
R4586 avdd.n82 avdd.n81 11.9049
R4587 avdd.n84 avdd.n83 11.9049
R4588 avdd.n71 avdd.n70 11.9049
R4589 avdd.n73 avdd.n72 11.9049
R4590 avdd.n60 avdd.n59 11.9049
R4591 avdd.n62 avdd.n61 11.9049
R4592 avdd.n49 avdd.n48 11.9049
R4593 avdd.n51 avdd.n50 11.9049
R4594 avdd.n38 avdd.n37 11.9049
R4595 avdd.n40 avdd.n39 11.9049
R4596 avdd.n27 avdd.n26 11.9049
R4597 avdd.n29 avdd.n28 11.9049
R4598 avdd.n16 avdd.n15 11.9049
R4599 avdd.n18 avdd.n17 11.9049
R4600 avdd.n5 avdd.n4 11.9049
R4601 avdd.n7 avdd.n6 11.9049
R4602 avdd.n170 avdd.n169 11.9049
R4603 avdd.n172 avdd.n171 11.9049
R4604 avdd.n159 avdd.n158 11.9049
R4605 avdd.n161 avdd.n160 11.9049
R4606 avdd.n148 avdd.n147 11.9049
R4607 avdd.n150 avdd.n149 11.9049
R4608 avdd.n137 avdd.n136 11.9049
R4609 avdd.n139 avdd.n138 11.9049
R4610 avdd.n126 avdd.n125 11.9049
R4611 avdd.n128 avdd.n127 11.9049
R4612 avdd.n115 avdd.n114 11.9049
R4613 avdd.n117 avdd.n116 11.9049
R4614 avdd.n104 avdd.n103 11.9049
R4615 avdd.n106 avdd.n105 11.9049
R4616 avdd.n93 avdd.n92 11.9049
R4617 avdd.n95 avdd.n94 11.9049
R4618 avdd.n258 avdd.n257 11.9049
R4619 avdd.n260 avdd.n259 11.9049
R4620 avdd.n247 avdd.n246 11.9049
R4621 avdd.n249 avdd.n248 11.9049
R4622 avdd.n236 avdd.n235 11.9049
R4623 avdd.n238 avdd.n237 11.9049
R4624 avdd.n225 avdd.n224 11.9049
R4625 avdd.n227 avdd.n226 11.9049
R4626 avdd.n214 avdd.n213 11.9049
R4627 avdd.n216 avdd.n215 11.9049
R4628 avdd.n203 avdd.n202 11.9049
R4629 avdd.n205 avdd.n204 11.9049
R4630 avdd.n192 avdd.n191 11.9049
R4631 avdd.n194 avdd.n193 11.9049
R4632 avdd.n181 avdd.n180 11.9049
R4633 avdd.n183 avdd.n182 11.9049
R4634 avdd.n302 avdd.n301 11.9049
R4635 avdd.n304 avdd.n303 11.9049
R4636 avdd.n291 avdd.n290 11.9049
R4637 avdd.n293 avdd.n292 11.9049
R4638 avdd.n280 avdd.n279 11.9049
R4639 avdd.n282 avdd.n281 11.9049
R4640 avdd.n269 avdd.n268 11.9049
R4641 avdd.n271 avdd.n270 11.9049
R4642 avdd.n407 avdd.t28 10.7165
R4643 avdd.n403 avdd.n402 6.48548
R4644 avdd.n403 avdd 4.8561
R4645 avdd.n83 avdd.t0 4.77693
R4646 avdd.t0 avdd.n82 4.77693
R4647 avdd.n72 avdd.t15 4.77693
R4648 avdd.t15 avdd.n71 4.77693
R4649 avdd.n61 avdd.t10 4.77693
R4650 avdd.t10 avdd.n60 4.77693
R4651 avdd.n50 avdd.t33 4.77693
R4652 avdd.t33 avdd.n49 4.77693
R4653 avdd.n39 avdd.t35 4.77693
R4654 avdd.t35 avdd.n38 4.77693
R4655 avdd.n28 avdd.t7 4.77693
R4656 avdd.t7 avdd.n27 4.77693
R4657 avdd.n17 avdd.t16 4.77693
R4658 avdd.t16 avdd.n16 4.77693
R4659 avdd.n6 avdd.t5 4.77693
R4660 avdd.t5 avdd.n5 4.77693
R4661 avdd.n171 avdd.t8 4.77693
R4662 avdd.t8 avdd.n170 4.77693
R4663 avdd.n160 avdd.t17 4.77693
R4664 avdd.t17 avdd.n159 4.77693
R4665 avdd.n149 avdd.t34 4.77693
R4666 avdd.t34 avdd.n148 4.77693
R4667 avdd.n138 avdd.t4 4.77693
R4668 avdd.t4 avdd.n137 4.77693
R4669 avdd.n127 avdd.t6 4.77693
R4670 avdd.t6 avdd.n126 4.77693
R4671 avdd.n116 avdd.t12 4.77693
R4672 avdd.t12 avdd.n115 4.77693
R4673 avdd.n105 avdd.t9 4.77693
R4674 avdd.t9 avdd.n104 4.77693
R4675 avdd.n94 avdd.t26 4.77693
R4676 avdd.t26 avdd.n93 4.77693
R4677 avdd.n259 avdd.t21 4.77693
R4678 avdd.t21 avdd.n258 4.77693
R4679 avdd.n248 avdd.t37 4.77693
R4680 avdd.t37 avdd.n247 4.77693
R4681 avdd.n237 avdd.t20 4.77693
R4682 avdd.t20 avdd.n236 4.77693
R4683 avdd.n226 avdd.t36 4.77693
R4684 avdd.t36 avdd.n225 4.77693
R4685 avdd.n215 avdd.t23 4.77693
R4686 avdd.t23 avdd.n214 4.77693
R4687 avdd.n204 avdd.t40 4.77693
R4688 avdd.t40 avdd.n203 4.77693
R4689 avdd.n193 avdd.t22 4.77693
R4690 avdd.t22 avdd.n192 4.77693
R4691 avdd.n182 avdd.t38 4.77693
R4692 avdd.t38 avdd.n181 4.77693
R4693 avdd.n303 avdd.t30 4.77693
R4694 avdd.t30 avdd.n302 4.77693
R4695 avdd.n292 avdd.t11 4.77693
R4696 avdd.t11 avdd.n291 4.77693
R4697 avdd.n281 avdd.t31 4.77693
R4698 avdd.t31 avdd.n280 4.77693
R4699 avdd.n270 avdd.t3 4.77693
R4700 avdd.t3 avdd.n269 4.77693
R4701 avdd.n406 avdd 3.12119
R4702 avdd.n405 avdd 3.12119
R4703 avdd.n404 avdd 3.12119
R4704 avdd avdd.n296 2.22787
R4705 avdd avdd.n274 2.22787
R4706 avdd.n10 avdd.n9 1.5505
R4707 avdd.n21 avdd.n20 1.5505
R4708 avdd.n32 avdd.n31 1.5505
R4709 avdd.n43 avdd.n42 1.5505
R4710 avdd.n54 avdd.n53 1.5505
R4711 avdd.n65 avdd.n64 1.5505
R4712 avdd.n76 avdd.n75 1.5505
R4713 avdd.n87 avdd.n86 1.5505
R4714 avdd.n98 avdd.n97 1.5505
R4715 avdd.n109 avdd.n108 1.5505
R4716 avdd.n120 avdd.n119 1.5505
R4717 avdd.n131 avdd.n130 1.5505
R4718 avdd.n142 avdd.n141 1.5505
R4719 avdd.n153 avdd.n152 1.5505
R4720 avdd.n164 avdd.n163 1.5505
R4721 avdd.n175 avdd.n174 1.5505
R4722 avdd.n186 avdd.n185 1.5505
R4723 avdd.n197 avdd.n196 1.5505
R4724 avdd.n208 avdd.n207 1.5505
R4725 avdd.n219 avdd.n218 1.5505
R4726 avdd.n230 avdd.n229 1.5505
R4727 avdd.n241 avdd.n240 1.5505
R4728 avdd.n252 avdd.n251 1.5505
R4729 avdd.n263 avdd.n262 1.5505
R4730 avdd.n274 avdd.n273 1.5505
R4731 avdd.n285 avdd.n284 1.5505
R4732 avdd.n296 avdd.n295 1.5505
R4733 avdd.n307 avdd.n306 1.5505
R4734 avdd.n354 avdd 1.38748
R4735 avdd.n378 avdd.n354 1.25871
R4736 avdd.n402 avdd.n378 1.25871
R4737 avdd.n87 avdd 1.24296
R4738 avdd.n76 avdd 1.24296
R4739 avdd.n65 avdd 1.24296
R4740 avdd.n54 avdd 1.24296
R4741 avdd.n43 avdd 1.24296
R4742 avdd.n32 avdd 1.24296
R4743 avdd.n21 avdd 1.24296
R4744 avdd.n10 avdd 1.24296
R4745 avdd.n175 avdd 1.24296
R4746 avdd.n164 avdd 1.24296
R4747 avdd.n153 avdd 1.24296
R4748 avdd.n142 avdd 1.24296
R4749 avdd.n131 avdd 1.24296
R4750 avdd.n120 avdd 1.24296
R4751 avdd.n109 avdd 1.24296
R4752 avdd.n98 avdd 1.24296
R4753 avdd.n263 avdd 1.24296
R4754 avdd.n252 avdd 1.24296
R4755 avdd.n241 avdd 1.24296
R4756 avdd.n230 avdd 1.24296
R4757 avdd.n219 avdd 1.24296
R4758 avdd.n208 avdd 1.24296
R4759 avdd.n197 avdd 1.24296
R4760 avdd.n186 avdd 1.24296
R4761 avdd.n307 avdd 1.24296
R4762 avdd.n296 avdd 1.24296
R4763 avdd.n285 avdd 1.24296
R4764 avdd.n274 avdd 1.24296
R4765 avdd avdd.n408 1.09544
R4766 avdd.n330 avdd.n329 0.645538
R4767 avdd.n353 avdd.n352 0.645538
R4768 avdd.n377 avdd.n376 0.645538
R4769 avdd.n401 avdd.n400 0.645538
R4770 avdd avdd.n87 0.492957
R4771 avdd avdd.n76 0.492957
R4772 avdd avdd.n65 0.492957
R4773 avdd avdd.n54 0.492957
R4774 avdd avdd.n43 0.492957
R4775 avdd avdd.n32 0.492957
R4776 avdd avdd.n21 0.492957
R4777 avdd avdd.n10 0.492957
R4778 avdd avdd.n175 0.492957
R4779 avdd avdd.n164 0.492957
R4780 avdd avdd.n153 0.492957
R4781 avdd avdd.n142 0.492957
R4782 avdd avdd.n131 0.492957
R4783 avdd avdd.n120 0.492957
R4784 avdd avdd.n109 0.492957
R4785 avdd avdd.n98 0.492957
R4786 avdd avdd.n263 0.492957
R4787 avdd avdd.n252 0.492957
R4788 avdd avdd.n241 0.492957
R4789 avdd avdd.n230 0.492957
R4790 avdd avdd.n219 0.492957
R4791 avdd avdd.n208 0.492957
R4792 avdd avdd.n197 0.492957
R4793 avdd avdd.n186 0.492957
R4794 avdd avdd.n307 0.492957
R4795 avdd avdd.n285 0.492957
R4796 avdd.n408 avdd.n407 0.426002
R4797 avdd.n408 avdd.n406 0.268357
R4798 avdd.n330 avdd.n308 0.265121
R4799 avdd.n353 avdd.n331 0.265121
R4800 avdd.n377 avdd.n355 0.265121
R4801 avdd.n401 avdd.n379 0.265121
R4802 avdd.n405 avdd.n404 0.148838
R4803 avdd.n404 avdd.n403 0.147954
R4804 avdd.n406 avdd.n405 0.144948
R4805 avdd.n354 avdd 0.129288
R4806 avdd.n378 avdd 0.128641
R4807 avdd.n402 avdd 0.128641
R4808 avdd.n329 avdd.n328 0.0554356
R4809 avdd.n352 avdd.n351 0.0554356
R4810 avdd.n376 avdd.n375 0.0554356
R4811 avdd.n400 avdd.n399 0.0554356
R4812 avdd avdd.n330 0.045098
R4813 avdd avdd.n353 0.045098
R4814 avdd avdd.n377 0.045098
R4815 avdd avdd.n401 0.045098
R4816 avdd.n407 avdd 0.0350686
R4817 multiplexer_0.vtrip_0.n0 multiplexer_0.vtrip_0.t1 41.2565
R4818 multiplexer_0.vtrip_0.n1 multiplexer_0.vtrip_0.n0 5.29988
R4819 multiplexer_0.vtrip_0.n1 multiplexer_0.vtrip_0.t6 16.8956
R4820 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n24 19.5921
R4821 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n1 1.62926
R4822 multiplexer_0.vtrip_0.n2 multiplexer_0.vtrip_0.n6 2.2505
R4823 multiplexer_0.vtrip_0.n7 multiplexer_0.vtrip_0.n11 2.2505
R4824 multiplexer_0.vtrip_0.n12 multiplexer_0.vtrip_0.n16 2.2505
R4825 multiplexer_0.vtrip_0.n2 multiplexer_0.vtrip_0.n23 2.85792
R4826 multiplexer_0.vtrip_0.n7 multiplexer_0.vtrip_0.n2 3.14503
R4827 multiplexer_0.vtrip_0.n24 multiplexer_0.vtrip_0.n7 2.97413
R4828 multiplexer_0.vtrip_0.n24 multiplexer_0.vtrip_0.n12 0.171398
R4829 multiplexer_0.vtrip_0.n12 multiplexer_0.vtrip_0.n20 2.84816
R4830 multiplexer_0.vtrip_0.n23 multiplexer_0.vtrip_0.t8 97.2843
R4831 multiplexer_0.vtrip_0.n23 multiplexer_0.vtrip_0.n22 2.41261
R4832 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n21 0.179071
R4833 multiplexer_0.vtrip_0.n22 multiplexer_0.vtrip_0.n21 1.66836
R4834 multiplexer_0.vtrip_0.n22 multiplexer_0.vtrip_0 1.07193
R4835 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.t7 18.1873
R4836 multiplexer_0.vtrip_0.n21 multiplexer_0.vtrip_0.t13 18.0088
R4837 multiplexer_0.vtrip_0.n20 multiplexer_0.vtrip_0.t14 97.2843
R4838 multiplexer_0.vtrip_0.n17 multiplexer_0.vtrip_0.n19 2.2505
R4839 multiplexer_0.vtrip_0.n20 multiplexer_0.vtrip_0.n17 0.172375
R4840 multiplexer_0.vtrip_0.n17 multiplexer_0.vtrip_0 0.103039
R4841 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n18 0.179071
R4842 multiplexer_0.vtrip_0.n19 multiplexer_0.vtrip_0.n18 1.66836
R4843 multiplexer_0.vtrip_0.n19 multiplexer_0.vtrip_0 1.07193
R4844 multiplexer_0.vtrip_0.t3 multiplexer_0.vtrip_0 18.5516
R4845 multiplexer_0.vtrip_0.n18 multiplexer_0.vtrip_0.t10 18.3731
R4846 multiplexer_0.vtrip_0.n14 multiplexer_0.vtrip_0.n13 1.5005
R4847 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n14 0.179071
R4848 multiplexer_0.vtrip_0.n16 multiplexer_0.vtrip_0.n14 1.66836
R4849 multiplexer_0.vtrip_0.n16 multiplexer_0.vtrip_0 1.07193
R4850 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n15 1.67907
R4851 multiplexer_0.vtrip_0.t18 multiplexer_0.vtrip_0.n15 16.8731
R4852 multiplexer_0.vtrip_0.n15 multiplexer_0.vtrip_0.t15 16.5088
R4853 multiplexer_0.vtrip_0.n13 multiplexer_0.vtrip_0.t9 16.8731
R4854 multiplexer_0.vtrip_0.n13 multiplexer_0.vtrip_0.t20 16.5088
R4855 multiplexer_0.vtrip_0.n9 multiplexer_0.vtrip_0.n8 1.5005
R4856 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n9 0.179071
R4857 multiplexer_0.vtrip_0.n11 multiplexer_0.vtrip_0.n9 1.66836
R4858 multiplexer_0.vtrip_0.n11 multiplexer_0.vtrip_0 1.07193
R4859 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n10 1.67907
R4860 multiplexer_0.vtrip_0.t12 multiplexer_0.vtrip_0.n10 16.8731
R4861 multiplexer_0.vtrip_0.n10 multiplexer_0.vtrip_0.t16 16.5088
R4862 multiplexer_0.vtrip_0.n8 multiplexer_0.vtrip_0.t19 16.8731
R4863 multiplexer_0.vtrip_0.n8 multiplexer_0.vtrip_0.t4 16.5088
R4864 multiplexer_0.vtrip_0.n4 multiplexer_0.vtrip_0.n3 1.5005
R4865 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n4 0.179071
R4866 multiplexer_0.vtrip_0.n6 multiplexer_0.vtrip_0.n4 1.66836
R4867 multiplexer_0.vtrip_0.n6 multiplexer_0.vtrip_0 1.07193
R4868 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0.n5 1.67907
R4869 multiplexer_0.vtrip_0.t17 multiplexer_0.vtrip_0.n5 16.8731
R4870 multiplexer_0.vtrip_0.n5 multiplexer_0.vtrip_0.t2 16.5088
R4871 multiplexer_0.vtrip_0.n3 multiplexer_0.vtrip_0.t5 16.8731
R4872 multiplexer_0.vtrip_0.n3 multiplexer_0.vtrip_0.t11 16.5088
R4873 multiplexer_0.vtrip_0.n0 multiplexer_0.vtrip_0.t0 227.385
R4874 multiplexer_0.in_1011.n0 multiplexer_0.in_1011.t2 228.216
R4875 multiplexer_0.in_1011.n0 multiplexer_0.in_1011.t0 83.695
R4876 multiplexer_0.in_1011.n3 multiplexer_0.in_1011.t1 10.5295
R4877 multiplexer_0.in_1011.n3 multiplexer_0.in_1011.t3 10.5285
R4878 multiplexer_0.in_1011.n2 multiplexer_0.in_1011.n1 4.33622
R4879 multiplexer_0.in_1011.n1 multiplexer_0.in_1011.n0 1.5005
R4880 multiplexer_0.in_1011 multiplexer_0.in_1011.n3 0.872792
R4881 multiplexer_0.in_1011.n1 multiplexer_0.in_1011 0.104667
R4882 multiplexer_0.in_1011.n2 multiplexer_0.in_1011 0.0166275
R4883 multiplexer_0.in_1011 multiplexer_0.in_1011.n2 0.00984659
R4884 multiplexer_0.trans_gate_m_21.in.t1 multiplexer_0.trans_gate_m_21.in.n0 228.216
R4885 multiplexer_0.trans_gate_m_21.in.n5 multiplexer_0.trans_gate_m_21.in.n0 1.5005
R4886 multiplexer_0.trans_gate_m_21.in.n0 multiplexer_0.trans_gate_m_21.in.t4 83.695
R4887 multiplexer_0.trans_gate_m_21.in multiplexer_0.trans_gate_m_21.in.n5 0.104667
R4888 multiplexer_0.trans_gate_m_21.in.n5 multiplexer_0.trans_gate_m_21.in.n4 4.43682
R4889 multiplexer_0.trans_gate_m_21.in.n2 multiplexer_0.trans_gate_m_21.in.n1 1.5005
R4890 multiplexer_0.trans_gate_m_21.in multiplexer_0.trans_gate_m_21.in.n2 0.104667
R4891 multiplexer_0.trans_gate_m_21.in.n4 multiplexer_0.trans_gate_m_21.in.n2 0.459875
R4892 multiplexer_0.trans_gate_m_21.in.n4 multiplexer_0.trans_gate_m_21.in 0.564042
R4893 multiplexer_0.trans_gate_m_21.in multiplexer_0.trans_gate_m_21.in.n3 1.60467
R4894 multiplexer_0.trans_gate_m_21.in.n3 multiplexer_0.trans_gate_m_21.in.t3 83.695
R4895 multiplexer_0.trans_gate_m_21.in.n3 multiplexer_0.trans_gate_m_21.in.t5 228.216
R4896 multiplexer_0.trans_gate_m_21.in.n1 multiplexer_0.trans_gate_m_21.in.t0 83.695
R4897 multiplexer_0.trans_gate_m_21.in.n1 multiplexer_0.trans_gate_m_21.in.t2 228.216
R4898 vtrip[1].n2 vtrip[1].t2 99.4021
R4899 vtrip[1].n0 vtrip[1].t0 23.1698
R4900 vtrip[1].n1 vtrip[1].t3 17.7681
R4901 vtrip[1].n0 vtrip[1].t1 17.7475
R4902 vtrip[1].n2 vtrip[1] 5.43617
R4903 vtrip[1].n3 vtrip[1].n2 1.7055
R4904 vtrip[1].n1 vtrip[1].n0 0.572059
R4905 vtrip[1].n3 vtrip[1].n1 0.1139
R4906 vtrip[1] vtrip[1].n3 0.0378665
R4907 comp_hyst_0.net5.n0 comp_hyst_0.net5.t2 44.0933
R4908 comp_hyst_0.net5.n7 comp_hyst_0.net5.n0 0.069579
R4909 comp_hyst_0.net5 comp_hyst_0.net5.n7 0.0436818
R4910 comp_hyst_0.net5.n2 comp_hyst_0.net5.n6 1.7055
R4911 comp_hyst_0.net5.n7 comp_hyst_0.net5.n2 0.751158
R4912 comp_hyst_0.net5.n2 comp_hyst_0.net5.n1 3.78196
R4913 comp_hyst_0.net5.n6 comp_hyst_0.net5.t5 5.24389
R4914 comp_hyst_0.net5.n6 comp_hyst_0.net5.n5 0.0929068
R4915 comp_hyst_0.net5.n5 comp_hyst_0.net5 0.0533418
R4916 comp_hyst_0.net5.n5 comp_hyst_0.net5.n3 5.69301
R4917 comp_hyst_0.net5.n4 comp_hyst_0.net5.n3 3.95781
R4918 comp_hyst_0.net5.n1 comp_hyst_0.net5.n4 3.95781
R4919 comp_hyst_0.net5.n1 comp_hyst_0.net5.t0 4.65803
R4920 comp_hyst_0.net5.t0 comp_hyst_0.net5.n3 4.65803
R4921 comp_hyst_0.net5.n4 comp_hyst_0.net5.t1 83.7172
R4922 comp_hyst_0.net5 comp_hyst_0.net5.t3 91.2731
R4923 comp_hyst_0.net5.n0 comp_hyst_0.net5.t4 87.9836
R4924 comp_hyst_0.net1.t1 comp_hyst_0.net1.n3 77.4826
R4925 comp_hyst_0.net1.n1 comp_hyst_0.net1.n3 1.46608
R4926 comp_hyst_0.net1.n2 comp_hyst_0.net1.n1 16.0859
R4927 comp_hyst_0.net1 comp_hyst_0.net1.n2 0.0178158
R4928 comp_hyst_0.net1.n2 comp_hyst_0.net1.t0 87.0947
R4929 comp_hyst_0.net1 comp_hyst_0.net1.n2 0.0247121
R4930 comp_hyst_0.net1 comp_hyst_0.net1.n2 0.0788333
R4931 comp_hyst_0.net1.n1 comp_hyst_0.net1.t3 77.4826
R4932 comp_hyst_0.net1.n3 comp_hyst_0.net1.n0 1.46608
R4933 comp_hyst_0.net1.n0 comp_hyst_0.net1.t4 78.9481
R4934 comp_hyst_0.net1.n0 comp_hyst_0.net1.t2 77.4826
R4935 multiplexer_0.in_0010.n0 multiplexer_0.in_0010.t0 228.216
R4936 multiplexer_0.in_0010.n0 multiplexer_0.in_0010.t2 83.695
R4937 multiplexer_0.in_0010.n4 multiplexer_0.in_0010.t1 10.5295
R4938 multiplexer_0.in_0010.n4 multiplexer_0.in_0010.t3 10.5285
R4939 multiplexer_0.in_0010 multiplexer_0.in_0010.n3 4.90529
R4940 multiplexer_0.in_0010.n2 multiplexer_0.in_0010.n1 4.34635
R4941 multiplexer_0.in_0010.n1 multiplexer_0.in_0010.n0 1.5005
R4942 multiplexer_0.in_0010 multiplexer_0.in_0010.n4 0.872792
R4943 multiplexer_0.in_0010.n3 multiplexer_0.in_0010 0.177654
R4944 multiplexer_0.in_0010.n1 multiplexer_0.in_0010 0.104667
R4945 multiplexer_0.in_0010.n2 multiplexer_0.in_0010 0.0064902
R4946 multiplexer_0.in_0010.n3 multiplexer_0.in_0010.n2 0.00411538
R4947 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t1 41.0738
R4948 multiplexer_0.vtrip_0_b.n1 multiplexer_0.vtrip_0_b.n0 4.08093
R4949 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n25 0.521333
R4950 multiplexer_0.vtrip_0_b.n25 multiplexer_0.vtrip_0_b.n1 2.87169
R4951 multiplexer_0.vtrip_0_b.n25 multiplexer_0.vtrip_0_b.t14 33.8377
R4952 multiplexer_0.vtrip_0_b.t14 multiplexer_0.vtrip_0_b.n24 33.8377
R4953 multiplexer_0.vtrip_0_b.n24 multiplexer_0.vtrip_0_b.n23 19.5721
R4954 multiplexer_0.vtrip_0_b.n1 multiplexer_0.vtrip_0_b.n24 2.69901
R4955 multiplexer_0.vtrip_0_b.n6 multiplexer_0.vtrip_0_b.n5 1.7055
R4956 multiplexer_0.vtrip_0_b.n11 multiplexer_0.vtrip_0_b.n10 1.7055
R4957 multiplexer_0.vtrip_0_b.n16 multiplexer_0.vtrip_0_b.n15 1.7055
R4958 multiplexer_0.vtrip_0_b.n21 multiplexer_0.vtrip_0_b.n20 1.7055
R4959 multiplexer_0.vtrip_0_b.n16 multiplexer_0.vtrip_0_b.n21 1.02307
R4960 multiplexer_0.vtrip_0_b.n11 multiplexer_0.vtrip_0_b.n16 1.02307
R4961 multiplexer_0.vtrip_0_b.n23 multiplexer_0.vtrip_0_b.n11 0.307905
R4962 multiplexer_0.vtrip_0_b.n23 multiplexer_0.vtrip_0_b.n6 0.715662
R4963 multiplexer_0.vtrip_0_b.n6 multiplexer_0.vtrip_0_b.n22 0.312351
R4964 multiplexer_0.vtrip_0_b.n21 multiplexer_0.vtrip_0_b.t2 99.4906
R4965 multiplexer_0.vtrip_0_b.n22 multiplexer_0.vtrip_0_b.t17 99.1756
R4966 multiplexer_0.vtrip_0_b.n22 multiplexer_0.vtrip_0_b 0.161507
R4967 multiplexer_0.vtrip_0_b.n18 multiplexer_0.vtrip_0_b.n17 1.5005
R4968 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n18 0.179071
R4969 multiplexer_0.vtrip_0_b.n20 multiplexer_0.vtrip_0_b.n18 1.66836
R4970 multiplexer_0.vtrip_0_b.n20 multiplexer_0.vtrip_0_b 1.07193
R4971 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n19 1.67907
R4972 multiplexer_0.vtrip_0_b.t19 multiplexer_0.vtrip_0_b.n19 16.8731
R4973 multiplexer_0.vtrip_0_b.n19 multiplexer_0.vtrip_0_b.t4 16.5088
R4974 multiplexer_0.vtrip_0_b.n17 multiplexer_0.vtrip_0_b.t8 16.8731
R4975 multiplexer_0.vtrip_0_b.n17 multiplexer_0.vtrip_0_b.t13 16.5088
R4976 multiplexer_0.vtrip_0_b.n13 multiplexer_0.vtrip_0_b.n12 1.5005
R4977 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n13 0.179071
R4978 multiplexer_0.vtrip_0_b.n15 multiplexer_0.vtrip_0_b.n13 1.66836
R4979 multiplexer_0.vtrip_0_b.n15 multiplexer_0.vtrip_0_b 1.07193
R4980 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n14 1.67907
R4981 multiplexer_0.vtrip_0_b.t12 multiplexer_0.vtrip_0_b.n14 16.8731
R4982 multiplexer_0.vtrip_0_b.n14 multiplexer_0.vtrip_0_b.t18 16.5088
R4983 multiplexer_0.vtrip_0_b.n12 multiplexer_0.vtrip_0_b.t3 16.8731
R4984 multiplexer_0.vtrip_0_b.n12 multiplexer_0.vtrip_0_b.t7 16.5088
R4985 multiplexer_0.vtrip_0_b.n8 multiplexer_0.vtrip_0_b.n7 1.5005
R4986 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n8 0.179071
R4987 multiplexer_0.vtrip_0_b.n10 multiplexer_0.vtrip_0_b.n8 1.66836
R4988 multiplexer_0.vtrip_0_b.n10 multiplexer_0.vtrip_0_b 1.07193
R4989 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n9 1.67907
R4990 multiplexer_0.vtrip_0_b.t6 multiplexer_0.vtrip_0_b.n9 16.8731
R4991 multiplexer_0.vtrip_0_b.n9 multiplexer_0.vtrip_0_b.t11 16.5088
R4992 multiplexer_0.vtrip_0_b.n7 multiplexer_0.vtrip_0_b.t15 16.8731
R4993 multiplexer_0.vtrip_0_b.n7 multiplexer_0.vtrip_0_b.t20 16.5088
R4994 multiplexer_0.vtrip_0_b.n3 multiplexer_0.vtrip_0_b.n2 1.5005
R4995 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n3 0.179071
R4996 multiplexer_0.vtrip_0_b.n5 multiplexer_0.vtrip_0_b.n3 1.66836
R4997 multiplexer_0.vtrip_0_b.n5 multiplexer_0.vtrip_0_b 1.07193
R4998 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_0_b.n4 1.67907
R4999 multiplexer_0.vtrip_0_b.t5 multiplexer_0.vtrip_0_b.n4 16.8731
R5000 multiplexer_0.vtrip_0_b.n4 multiplexer_0.vtrip_0_b.t9 16.5088
R5001 multiplexer_0.vtrip_0_b.n2 multiplexer_0.vtrip_0_b.t10 16.8731
R5002 multiplexer_0.vtrip_0_b.n2 multiplexer_0.vtrip_0_b.t16 16.5088
R5003 multiplexer_0.vtrip_0_b.n0 multiplexer_0.vtrip_0_b.t0 227.512
R5004 a_n12118_2955.t0 a_n12118_2955.t1 21.2567
R5005 a_n8898_3333.t0 a_n8898_3333.t1 21.167
R5006 voltage_divider_0.51.n0 voltage_divider_0.51.t0 10.6833
R5007 voltage_divider_0.51.n0 voltage_divider_0.51.t1 10.5739
R5008 voltage_divider_0.51 voltage_divider_0.51.n0 0.036669
R5009 multiplexer_0.in_0000.n0 multiplexer_0.in_0000.t0 228.216
R5010 multiplexer_0.in_0000.n0 multiplexer_0.in_0000.t3 83.695
R5011 multiplexer_0.in_0000.n3 multiplexer_0.in_0000.t1 10.5295
R5012 multiplexer_0.in_0000.n3 multiplexer_0.in_0000.t2 10.5285
R5013 multiplexer_0.in_0000 multiplexer_0.in_0000.n2 5.93817
R5014 multiplexer_0.in_0000 multiplexer_0.in_0000.n0 1.60467
R5015 multiplexer_0.in_0000 multiplexer_0.in_0000.n3 0.872792
R5016 multiplexer_0.in_0000.n2 multiplexer_0.in_0000 0.471654
R5017 multiplexer_0.in_0000.n1 multiplexer_0.in_0000 0.414042
R5018 multiplexer_0.in_0000.n1 multiplexer_0.in_0000 0.0140417
R5019 multiplexer_0.in_0000.n2 multiplexer_0.in_0000.n1 0.0101154
R5020 vin.t0 vin.n0 228.216
R5021 vin.n7 vin.n0 1.5005
R5022 vin.n0 vin.t2 83.695
R5023 vin vin.n7 0.104667
R5024 vin.n7 vin.n1 2.26752
R5025 vin.n1 vin 0.156447
R5026 vin vin.n6 2.47322
R5027 vin.n5 vin.n6 1.5005
R5028 vin vin.n6 0.104667
R5029 vin.t3 vin.n5 83.695
R5030 vin.t1 vin.n5 228.216
R5031 vin.n1 vin 12.6632
R5032 vin vin.n4 11.7757
R5033 vin vin.n4 2.0685
R5034 vin vin.n4 0.00103107
R5035 vin.n4 vin.n2 0.0129802
R5036 vin.n2 vin.n3 0.475071
R5037 vin.t4 vin.n3 8.09606
R5038 vin.n3 vin.t5 8.26823
R5039 vin.t6 vin.n2 101.106
R5040 a_n15874_13161.t0 a_n15874_13161.t1 21.2567
R5041 a_n12654_13539.t0 a_n12654_13539.t1 21.167
R5042 multiplexer_0.in_1001.n0 multiplexer_0.in_1001.t3 228.216
R5043 multiplexer_0.in_1001.n0 multiplexer_0.in_1001.t0 83.695
R5044 multiplexer_0.in_1001.n2 multiplexer_0.in_1001.t1 10.5295
R5045 multiplexer_0.in_1001.n2 multiplexer_0.in_1001.t2 10.5285
R5046 multiplexer_0.in_1001 multiplexer_0.in_1001.n1 2.54596
R5047 multiplexer_0.in_1001 multiplexer_0.in_1001.n0 1.60467
R5048 multiplexer_0.in_1001 multiplexer_0.in_1001.n2 0.872792
R5049 multiplexer_0.in_1001.n1 multiplexer_0.in_1001 0.3505
R5050 multiplexer_0.in_1001.n1 multiplexer_0.in_1001 0.0775833
R5051 multiplexer_0.trans_gate_m_23.in.t1 multiplexer_0.trans_gate_m_23.in.n0 228.216
R5052 multiplexer_0.trans_gate_m_23.in.n6 multiplexer_0.trans_gate_m_23.in.n0 1.5005
R5053 multiplexer_0.trans_gate_m_23.in.n0 multiplexer_0.trans_gate_m_23.in.t4 83.695
R5054 multiplexer_0.trans_gate_m_23.in multiplexer_0.trans_gate_m_23.in.n6 0.104667
R5055 multiplexer_0.trans_gate_m_23.in.n3 multiplexer_0.trans_gate_m_23.in.n4 10.4956
R5056 multiplexer_0.trans_gate_m_23.in.n3 multiplexer_0.trans_gate_m_23.in.n2 2.45249
R5057 multiplexer_0.trans_gate_m_23.in.n6 multiplexer_0.trans_gate_m_23.in.n3 2.44157
R5058 multiplexer_0.trans_gate_m_23.in.n4 multiplexer_0.trans_gate_m_23.in.n5 1.5005
R5059 multiplexer_0.trans_gate_m_23.in multiplexer_0.trans_gate_m_23.in.n4 0.104667
R5060 multiplexer_0.trans_gate_m_23.in.n5 multiplexer_0.trans_gate_m_23.in.t5 83.695
R5061 multiplexer_0.trans_gate_m_23.in.n5 multiplexer_0.trans_gate_m_23.in.t2 228.216
R5062 multiplexer_0.trans_gate_m_23.in.n2 multiplexer_0.trans_gate_m_23.in.n1 1.5005
R5063 multiplexer_0.trans_gate_m_23.in multiplexer_0.trans_gate_m_23.in.n2 0.104667
R5064 multiplexer_0.trans_gate_m_23.in.n1 multiplexer_0.trans_gate_m_23.in.t0 83.695
R5065 multiplexer_0.trans_gate_m_23.in.n1 multiplexer_0.trans_gate_m_23.in.t3 228.216
R5066 a_n8362_13161.t0 a_n8362_13161.t1 21.2567
R5067 a_n5142_12783.t0 a_n5142_12783.t1 21.167
R5068 a_n12118_7491.t0 a_n12118_7491.t1 21.2567
R5069 a_n8898_7113.t0 a_n8898_7113.t1 21.167
R5070 multiplexer_0.vtrip_2_b.n0 multiplexer_0.vtrip_2_b.t0 41.0738
R5071 multiplexer_0.vtrip_2_b.n1 multiplexer_0.vtrip_2_b.n0 4.08093
R5072 multiplexer_0.vtrip_2_b multiplexer_0.vtrip_2_b.n8 0.521333
R5073 multiplexer_0.vtrip_2_b.n8 multiplexer_0.vtrip_2_b.n1 2.87169
R5074 multiplexer_0.vtrip_2_b.n8 multiplexer_0.vtrip_2_b.t2 33.8377
R5075 multiplexer_0.vtrip_2_b.t2 multiplexer_0.vtrip_2_b.n7 33.8377
R5076 multiplexer_0.vtrip_2_b.n7 multiplexer_0.vtrip_2_b.n6 13.7788
R5077 multiplexer_0.vtrip_2_b.n1 multiplexer_0.vtrip_2_b.n7 2.69901
R5078 multiplexer_0.vtrip_2_b.n6 multiplexer_0.vtrip_2_b.n2 0.456527
R5079 multiplexer_0.vtrip_2_b.n2 multiplexer_0.vtrip_2_b.n5 0.536237
R5080 multiplexer_0.vtrip_2_b.n5 multiplexer_0.vtrip_2_b.t6 99.1792
R5081 multiplexer_0.vtrip_2_b.n5 multiplexer_0.vtrip_2_b.n4 0.437791
R5082 multiplexer_0.vtrip_2_b.n4 multiplexer_0.vtrip_2_b.n3 0.511784
R5083 multiplexer_0.vtrip_2_b multiplexer_0.vtrip_2_b.n3 0.546399
R5084 multiplexer_0.vtrip_2_b.n4 multiplexer_0.vtrip_2_b 2.77693
R5085 multiplexer_0.vtrip_2_b.t7 multiplexer_0.vtrip_2_b 18.5516
R5086 multiplexer_0.vtrip_2_b.n3 multiplexer_0.vtrip_2_b 2.77693
R5087 multiplexer_0.vtrip_2_b multiplexer_0.vtrip_2_b.t5 18.1873
R5088 multiplexer_0.vtrip_2_b.n6 multiplexer_0.vtrip_2_b 2.83219
R5089 multiplexer_0.vtrip_2_b.t3 multiplexer_0.vtrip_2_b 18.5516
R5090 multiplexer_0.vtrip_2_b.n2 multiplexer_0.vtrip_2_b 2.77693
R5091 multiplexer_0.vtrip_2_b multiplexer_0.vtrip_2_b.t4 18.1873
R5092 multiplexer_0.vtrip_2_b.n0 multiplexer_0.vtrip_2_b.t1 227.512
R5093 a_n15874_3333.t0 a_n15874_3333.t1 21.2567
R5094 a_n12654_3711.t0 a_n12654_3711.t1 21.167
R5095 a_n8898_n447.t0 a_n8898_n447.t1 21.341
R5096 a_n5142_n825.t0 a_n5142_n825.t1 21.167
R5097 vbg.n1 vbg.t2 101.106
R5098 vbg.n0 vbg.t1 8.61346
R5099 vbg.n0 vbg.t0 8.09814
R5100 vbg.n2 vbg 4.75829
R5101 vbg vbg.n2 2.0685
R5102 vbg.n1 vbg.n0 0.303134
R5103 vbg.n2 vbg.n1 0.0129802
R5104 vbg.n2 vbg 0.00103107
R5105 a_n12118_10515.t0 a_n12118_10515.t1 21.2567
R5106 a_n8898_10893.t0 a_n8898_10893.t1 21.167
R5107 a_n8362_8625.t0 a_n8362_8625.t1 21.2567
R5108 multiplexer_0.in_0100.n0 multiplexer_0.in_0100.t1 228.216
R5109 multiplexer_0.in_0100.n0 multiplexer_0.in_0100.t3 83.695
R5110 multiplexer_0.in_0100.n3 multiplexer_0.in_0100.t2 10.5739
R5111 multiplexer_0.in_0100.n3 multiplexer_0.in_0100.t0 10.5739
R5112 multiplexer_0.in_0100 multiplexer_0.in_0100.n2 5.1017
R5113 multiplexer_0.in_0100 multiplexer_0.in_0100.n3 2.20538
R5114 multiplexer_0.in_0100 multiplexer_0.in_0100.n0 1.60467
R5115 multiplexer_0.in_0100.n2 multiplexer_0.in_0100 0.471654
R5116 multiplexer_0.in_0100.n1 multiplexer_0.in_0100 0.414042
R5117 multiplexer_0.in_0100.n1 multiplexer_0.in_0100 0.0140417
R5118 multiplexer_0.in_0100.n2 multiplexer_0.in_0100.n1 0.0101154
R5119 a_n5142_5979.t0 a_n5142_5979.t1 21.0576
R5120 a_n15874_10893.t0 a_n15874_10893.t1 21.2567
R5121 a_n12654_11271.t0 a_n12654_11271.t1 21.167
R5122 multiplexer_0.in_0101.n0 multiplexer_0.in_0101.t3 228.216
R5123 multiplexer_0.in_0101.n0 multiplexer_0.in_0101.t0 83.695
R5124 multiplexer_0.in_0101.n3 multiplexer_0.in_0101.t2 10.5739
R5125 multiplexer_0.in_0101.n3 multiplexer_0.in_0101.t1 10.5739
R5126 multiplexer_0.in_0101 multiplexer_0.in_0101.n2 4.09284
R5127 multiplexer_0.in_0101 multiplexer_0.in_0101.n3 2.20538
R5128 multiplexer_0.in_0101 multiplexer_0.in_0101.n0 1.60467
R5129 multiplexer_0.in_0101.n2 multiplexer_0.in_0101 0.471654
R5130 multiplexer_0.in_0101.n1 multiplexer_0.in_0101 0.414042
R5131 multiplexer_0.in_0101.n1 multiplexer_0.in_0101 0.0140417
R5132 multiplexer_0.in_0101.n2 multiplexer_0.in_0101.n1 0.0101154
R5133 multiplexer_0.trans_gate_m_27.in.t0 multiplexer_0.trans_gate_m_27.in.n0 228.216
R5134 multiplexer_0.trans_gate_m_27.in.n6 multiplexer_0.trans_gate_m_27.in.n0 1.5005
R5135 multiplexer_0.trans_gate_m_27.in.n0 multiplexer_0.trans_gate_m_27.in.t3 83.695
R5136 multiplexer_0.trans_gate_m_27.in multiplexer_0.trans_gate_m_27.in.n6 0.104667
R5137 multiplexer_0.trans_gate_m_27.in.n3 multiplexer_0.trans_gate_m_27.in.n4 10.4956
R5138 multiplexer_0.trans_gate_m_27.in.n3 multiplexer_0.trans_gate_m_27.in.n2 2.45249
R5139 multiplexer_0.trans_gate_m_27.in.n6 multiplexer_0.trans_gate_m_27.in.n3 2.44157
R5140 multiplexer_0.trans_gate_m_27.in.n4 multiplexer_0.trans_gate_m_27.in.n5 1.5005
R5141 multiplexer_0.trans_gate_m_27.in multiplexer_0.trans_gate_m_27.in.n4 0.104667
R5142 multiplexer_0.trans_gate_m_27.in.n5 multiplexer_0.trans_gate_m_27.in.t5 83.695
R5143 multiplexer_0.trans_gate_m_27.in.n5 multiplexer_0.trans_gate_m_27.in.t2 228.216
R5144 multiplexer_0.trans_gate_m_27.in.n2 multiplexer_0.trans_gate_m_27.in.n1 1.5005
R5145 multiplexer_0.trans_gate_m_27.in multiplexer_0.trans_gate_m_27.in.n2 0.104667
R5146 multiplexer_0.trans_gate_m_27.in.n1 multiplexer_0.trans_gate_m_27.in.t1 83.695
R5147 multiplexer_0.trans_gate_m_27.in.n1 multiplexer_0.trans_gate_m_27.in.t4 228.216
R5148 a_n8362_10137.t0 a_n8362_10137.t1 21.2567
R5149 a_n5142_9759.t0 a_n5142_9759.t1 21.167
R5150 a_n12118_6735.t0 a_n12118_6735.t1 21.2567
R5151 multiplexer_0.trans_gate_m_28.in.n0 multiplexer_0.trans_gate_m_28.in.t0 228.216
R5152 multiplexer_0.trans_gate_m_28.in.n0 multiplexer_0.trans_gate_m_28.in.t3 83.695
R5153 multiplexer_0.trans_gate_m_28.in.n5 multiplexer_0.trans_gate_m_28.in.n4 1.5005
R5154 multiplexer_0.trans_gate_m_28.in multiplexer_0.trans_gate_m_28.in.n5 0.104667
R5155 multiplexer_0.trans_gate_m_28.in.n5 multiplexer_0.trans_gate_m_28.in.n3 0.459875
R5156 multiplexer_0.trans_gate_m_28.in.n3 multiplexer_0.trans_gate_m_28.in 0.553625
R5157 multiplexer_0.trans_gate_m_28.in multiplexer_0.trans_gate_m_28.in.n0 1.60467
R5158 multiplexer_0.trans_gate_m_28.in.n4 multiplexer_0.trans_gate_m_28.in.t1 83.695
R5159 multiplexer_0.trans_gate_m_28.in.n4 multiplexer_0.trans_gate_m_28.in.t4 228.216
R5160 multiplexer_0.trans_gate_m_28.in.n3 multiplexer_0.trans_gate_m_28.in.n2 4.43682
R5161 multiplexer_0.trans_gate_m_28.in.n2 multiplexer_0.trans_gate_m_28.in.n1 1.5005
R5162 multiplexer_0.trans_gate_m_28.in multiplexer_0.trans_gate_m_28.in.n2 0.104667
R5163 multiplexer_0.trans_gate_m_28.in.n1 multiplexer_0.trans_gate_m_28.in.t5 83.695
R5164 multiplexer_0.trans_gate_m_28.in.n1 multiplexer_0.trans_gate_m_28.in.t2 228.216
R5165 ena.n9 ena.t6 99.4005
R5166 ena.n11 ena.t2 99.4005
R5167 ena.n1 ena.t7 35.2949
R5168 ena.n2 ena.t7 35.2949
R5169 ena.t3 ena.n0 34.8146
R5170 ena.n3 ena.t3 34.8146
R5171 ena.n2 ena.t1 33.8377
R5172 ena.t1 ena.n1 33.8377
R5173 ena ena.t0 25.2266
R5174 ena.n8 ena.t5 20.4065
R5175 ena.n6 ena.t5 19.344
R5176 ena.n5 ena.t4 17.6981
R5177 ena.n11 ena.n10 9.6297
R5178 ena.n10 ena 3.99824
R5179 ena.n6 ena.n5 3.48479
R5180 ena.n7 ena.n6 2.7271
R5181 ena.n4 ena.n0 1.8089
R5182 ena.n4 ena.n3 1.7055
R5183 ena.n8 ena.n7 1.7055
R5184 ena.n1 ena.n0 1.07287
R5185 ena.n3 ena.n2 1.07287
R5186 ena.n10 ena 0.46101
R5187 ena.n9 ena.n8 0.373074
R5188 ena.n5 ena.n4 0.16323
R5189 ena ena.n11 0.063
R5190 ena ena.n9 0.0309688
R5191 ena.n7 ena 0.0115247
R5192 a_n5142_n1959.t1 a_n5142_n1959.t0 41.7607
R5193 a_n12118_4467.t0 a_n12118_4467.t1 21.2567
R5194 a_n8898_4089.t0 a_n8898_4089.t1 21.167
R5195 a_n15874_1065.t0 a_n15874_1065.t1 21.2567
R5196 a_n12654_1065.t0 a_n12654_1065.t1 21.341
R5197 multiplexer_0.vtrip_3_b.n0 multiplexer_0.vtrip_3_b.t1 41.0738
R5198 multiplexer_0.vtrip_3_b.n1 multiplexer_0.vtrip_3_b.n0 5.5069
R5199 multiplexer_0.vtrip_3_b multiplexer_0.vtrip_3_b.n1 1.82794
R5200 multiplexer_0.vtrip_3_b multiplexer_0.vtrip_3_b.n3 0.545128
R5201 multiplexer_0.vtrip_3_b.t4 multiplexer_0.vtrip_3_b.n3 99.2037
R5202 multiplexer_0.vtrip_3_b.n3 multiplexer_0.vtrip_3_b 2.77693
R5203 multiplexer_0.vtrip_3_b multiplexer_0.vtrip_3_b.n2 1.67907
R5204 multiplexer_0.vtrip_3_b.t5 multiplexer_0.vtrip_3_b.n2 16.8731
R5205 multiplexer_0.vtrip_3_b.n2 multiplexer_0.vtrip_3_b.t3 16.5088
R5206 multiplexer_0.vtrip_3_b.n1 multiplexer_0.vtrip_3_b.t2 16.8829
R5207 multiplexer_0.vtrip_3_b.n0 multiplexer_0.vtrip_3_b.t0 227.512
R5208 multiplexer_0.trans_gate_m_33.in.t0 multiplexer_0.trans_gate_m_33.in.n0 228.216
R5209 multiplexer_0.trans_gate_m_33.in.n5 multiplexer_0.trans_gate_m_33.in.n0 1.5005
R5210 multiplexer_0.trans_gate_m_33.in.n0 multiplexer_0.trans_gate_m_33.in.t4 83.695
R5211 multiplexer_0.trans_gate_m_33.in multiplexer_0.trans_gate_m_33.in.n5 0.104667
R5212 multiplexer_0.trans_gate_m_33.in.n5 multiplexer_0.trans_gate_m_33.in.n3 0.459875
R5213 multiplexer_0.trans_gate_m_33.in.n3 multiplexer_0.trans_gate_m_33.in 0.563
R5214 multiplexer_0.trans_gate_m_33.in multiplexer_0.trans_gate_m_33.in.n4 1.60467
R5215 multiplexer_0.trans_gate_m_33.in.n4 multiplexer_0.trans_gate_m_33.in.t2 83.695
R5216 multiplexer_0.trans_gate_m_33.in.n4 multiplexer_0.trans_gate_m_33.in.t3 228.216
R5217 multiplexer_0.trans_gate_m_33.in.n3 multiplexer_0.trans_gate_m_33.in.n2 5.41376
R5218 multiplexer_0.trans_gate_m_33.in.n2 multiplexer_0.trans_gate_m_33.in.n1 1.5005
R5219 multiplexer_0.trans_gate_m_33.in multiplexer_0.trans_gate_m_33.in.n2 0.104667
R5220 multiplexer_0.trans_gate_m_33.in.n1 multiplexer_0.trans_gate_m_33.in.t1 83.695
R5221 multiplexer_0.trans_gate_m_33.in.n1 multiplexer_0.trans_gate_m_33.in.t5 228.216
R5222 a_n8362_13917.t0 a_n8362_13917.t1 21.2567
R5223 a_n5142_14295.t0 a_n5142_14295.t1 21.167
R5224 a_n8898_10137.t0 a_n8898_10137.t1 21.167
R5225 a_n5142_13539.t0 a_n5142_13539.t1 21.167
R5226 multiplexer_0.in_1010.n0 multiplexer_0.in_1010.t0 228.216
R5227 multiplexer_0.in_1010.n0 multiplexer_0.in_1010.t3 83.695
R5228 multiplexer_0.in_1010.n4 multiplexer_0.in_1010.t2 10.5739
R5229 multiplexer_0.in_1010.n4 multiplexer_0.in_1010.t1 10.5739
R5230 multiplexer_0.in_1010.n2 multiplexer_0.in_1010.n1 4.34635
R5231 multiplexer_0.in_1010 multiplexer_0.in_1010.n3 3.97588
R5232 multiplexer_0.in_1010 multiplexer_0.in_1010.n4 2.20538
R5233 multiplexer_0.in_1010.n1 multiplexer_0.in_1010.n0 1.5005
R5234 multiplexer_0.in_1010.n3 multiplexer_0.in_1010 0.177654
R5235 multiplexer_0.in_1010.n1 multiplexer_0.in_1010 0.104667
R5236 multiplexer_0.in_1010.n2 multiplexer_0.in_1010 0.0064902
R5237 multiplexer_0.in_1010.n3 multiplexer_0.in_1010.n2 0.00411538
R5238 a_n12654_n69.t0 a_n12654_n69.t1 21.34
R5239 a_n15874_4845.t0 a_n15874_4845.t1 21.2567
R5240 a_n12654_4467.t0 a_n12654_4467.t1 21.167
R5241 comp_hyst_0.ena_b.n0 comp_hyst_0.ena_b.t1 83.7172
R5242 comp_hyst_0.ena_b comp_hyst_0.ena_b.n0 0.38198
R5243 comp_hyst_0.ena_b comp_hyst_0.ena_b.n9 0.0575652
R5244 comp_hyst_0.ena_b comp_hyst_0.ena_b.n9 0.137405
R5245 comp_hyst_0.ena_b.n9 comp_hyst_0.ena_b.n8 0.997524
R5246 comp_hyst_0.ena_b comp_hyst_0.ena_b.n8 0.314856
R5247 comp_hyst_0.ena_b.n8 comp_hyst_0.ena_b.t0 228.338
R5248 comp_hyst_0.ena_b.n2 comp_hyst_0.ena_b.n1 1.7055
R5249 comp_hyst_0.ena_b.n0 comp_hyst_0.ena_b.n2 3.37881
R5250 comp_hyst_0.ena_b.n2 comp_hyst_0.ena_b.n3 3.01285
R5251 comp_hyst_0.ena_b.n3 comp_hyst_0.ena_b.n4 1.45774
R5252 comp_hyst_0.ena_b.n4 comp_hyst_0.ena_b.t4 34.5866
R5253 comp_hyst_0.ena_b.n6 comp_hyst_0.ena_b.t4 34.5866
R5254 comp_hyst_0.ena_b.n1 comp_hyst_0.ena_b.n7 2.81589
R5255 comp_hyst_0.ena_b.n1 comp_hyst_0.ena_b.n5 1.20445
R5256 comp_hyst_0.ena_b.n5 comp_hyst_0.ena_b.n6 1.45774
R5257 comp_hyst_0.ena_b.n7 comp_hyst_0.ena_b 0.0481042
R5258 comp_hyst_0.ena_b.n7 comp_hyst_0.ena_b.t5 23.3374
R5259 comp_hyst_0.ena_b.n6 comp_hyst_0.ena_b.t3 33.1294
R5260 comp_hyst_0.ena_b.n4 comp_hyst_0.ena_b.t3 33.1294
R5261 comp_hyst_0.ena_b.n5 comp_hyst_0.ena_b.t2 33.1294
R5262 comp_hyst_0.ena_b.n3 comp_hyst_0.ena_b.t2 33.1294
R5263 a_n12118_14295.t0 a_n12118_14295.t1 21.2567
R5264 a_n8898_14673.t0 a_n8898_14673.t1 21.341
R5265 vtrip[2].n2 vtrip[2].t3 99.4021
R5266 vtrip[2].n0 vtrip[2].t2 23.1698
R5267 vtrip[2].n1 vtrip[2].t1 17.7681
R5268 vtrip[2].n0 vtrip[2].t0 17.7475
R5269 vtrip[2].n2 vtrip[2] 5.20458
R5270 vtrip[2].n3 vtrip[2].n2 1.7055
R5271 vtrip[2].n1 vtrip[2].n0 0.572059
R5272 vtrip[2].n3 vtrip[2].n1 0.1139
R5273 vtrip[2] vtrip[2].n3 0.0378665
R5274 level_shifter_2.in_b.n0 level_shifter_2.in_b.t1 83.7172
R5275 level_shifter_2.in_b.n0 level_shifter_2.in_b.t0 229.644
R5276 level_shifter_2.in_b level_shifter_2.in_b.n0 5.2032
R5277 level_shifter_2.in_b level_shifter_2.in_b.t2 21.9226
R5278 a_n12654_1821.t0 a_n12654_1821.t1 21.341
R5279 a_n8898_1821.t0 a_n8898_1821.t1 21.167
R5280 a_n15874_14673.t0 a_n15874_14673.t1 21.2567
R5281 a_n12654_15051.t0 a_n12654_15051.t1 21.34
R5282 multiplexer_0.trans_gate_m_18.in.t1 multiplexer_0.trans_gate_m_18.in.n0 228.216
R5283 multiplexer_0.trans_gate_m_18.in.n6 multiplexer_0.trans_gate_m_18.in.n0 1.5005
R5284 multiplexer_0.trans_gate_m_18.in.n0 multiplexer_0.trans_gate_m_18.in.t4 83.695
R5285 multiplexer_0.trans_gate_m_18.in multiplexer_0.trans_gate_m_18.in.n6 0.104667
R5286 multiplexer_0.trans_gate_m_18.in.n3 multiplexer_0.trans_gate_m_18.in.n4 10.4956
R5287 multiplexer_0.trans_gate_m_18.in.n3 multiplexer_0.trans_gate_m_18.in.n2 2.45249
R5288 multiplexer_0.trans_gate_m_18.in.n6 multiplexer_0.trans_gate_m_18.in.n3 2.44157
R5289 multiplexer_0.trans_gate_m_18.in.n4 multiplexer_0.trans_gate_m_18.in.n5 1.5005
R5290 multiplexer_0.trans_gate_m_18.in multiplexer_0.trans_gate_m_18.in.n4 0.104667
R5291 multiplexer_0.trans_gate_m_18.in.n5 multiplexer_0.trans_gate_m_18.in.t5 83.695
R5292 multiplexer_0.trans_gate_m_18.in.n5 multiplexer_0.trans_gate_m_18.in.t2 228.216
R5293 multiplexer_0.trans_gate_m_18.in.n2 multiplexer_0.trans_gate_m_18.in.n1 1.5005
R5294 multiplexer_0.trans_gate_m_18.in multiplexer_0.trans_gate_m_18.in.n2 0.104667
R5295 multiplexer_0.trans_gate_m_18.in.n1 multiplexer_0.trans_gate_m_18.in.t0 83.695
R5296 multiplexer_0.trans_gate_m_18.in.n1 multiplexer_0.trans_gate_m_18.in.t3 228.216
R5297 a_n12118_8247.t0 a_n12118_8247.t1 21.2567
R5298 a_n8898_7869.t0 a_n8898_7869.t1 21.167
R5299 multiplexer_0.in_1110.n0 multiplexer_0.in_1110.t0 228.216
R5300 multiplexer_0.in_1110.n0 multiplexer_0.in_1110.t3 83.695
R5301 multiplexer_0.in_1110.n4 multiplexer_0.in_1110.t2 10.5739
R5302 multiplexer_0.in_1110.n4 multiplexer_0.in_1110.t1 10.5739
R5303 multiplexer_0.in_1110.n2 multiplexer_0.in_1110.n1 4.34635
R5304 multiplexer_0.in_1110 multiplexer_0.in_1110.n3 3.28049
R5305 multiplexer_0.in_1110 multiplexer_0.in_1110.n4 2.20538
R5306 multiplexer_0.in_1110.n1 multiplexer_0.in_1110.n0 1.5005
R5307 multiplexer_0.in_1110.n3 multiplexer_0.in_1110 0.177654
R5308 multiplexer_0.in_1110.n1 multiplexer_0.in_1110 0.104667
R5309 multiplexer_0.in_1110.n2 multiplexer_0.in_1110 0.0064902
R5310 multiplexer_0.in_1110.n3 multiplexer_0.in_1110.n2 0.00411538
R5311 multiplexer_0.trans_gate_m_19.in.t0 multiplexer_0.trans_gate_m_19.in.n0 228.216
R5312 multiplexer_0.trans_gate_m_19.in.n5 multiplexer_0.trans_gate_m_19.in.n0 1.5005
R5313 multiplexer_0.trans_gate_m_19.in.n0 multiplexer_0.trans_gate_m_19.in.t3 83.695
R5314 multiplexer_0.trans_gate_m_19.in multiplexer_0.trans_gate_m_19.in.n5 0.104667
R5315 multiplexer_0.trans_gate_m_19.in.n5 multiplexer_0.trans_gate_m_19.in.n4 4.43682
R5316 multiplexer_0.trans_gate_m_19.in.n2 multiplexer_0.trans_gate_m_19.in.n1 1.5005
R5317 multiplexer_0.trans_gate_m_19.in multiplexer_0.trans_gate_m_19.in.n2 0.104667
R5318 multiplexer_0.trans_gate_m_19.in.n4 multiplexer_0.trans_gate_m_19.in.n2 0.459875
R5319 multiplexer_0.trans_gate_m_19.in.n4 multiplexer_0.trans_gate_m_19.in 0.564042
R5320 multiplexer_0.trans_gate_m_19.in multiplexer_0.trans_gate_m_19.in.n3 1.60467
R5321 multiplexer_0.trans_gate_m_19.in.n3 multiplexer_0.trans_gate_m_19.in.t2 83.695
R5322 multiplexer_0.trans_gate_m_19.in.n3 multiplexer_0.trans_gate_m_19.in.t5 228.216
R5323 multiplexer_0.trans_gate_m_19.in.n1 multiplexer_0.trans_gate_m_19.in.t1 83.695
R5324 multiplexer_0.trans_gate_m_19.in.n1 multiplexer_0.trans_gate_m_19.in.t4 228.216
R5325 comp_hyst_0.net2 comp_hyst_0.net2.t0 232.147
R5326 comp_hyst_0.net2 comp_hyst_0.net2.t1 90.5793
R5327 comp_hyst_0.net2 comp_hyst_0.net2.t2 86.8087
R5328 comp_hyst_0.net2 comp_hyst_0.net2.t3 84.6545
R5329 a_n15874_n1959.t0 a_n15874_n1959.t1 21.2567
R5330 a_n12654_n1959.t0 a_n12654_n1959.t1 21.341
R5331 a_n8898_1065.t0 a_n8898_1065.t1 21.34
R5332 a_n5142_687.t0 a_n5142_687.t1 21.167
R5333 multiplexer_0.in_0011.n0 multiplexer_0.in_0011.t3 228.216
R5334 multiplexer_0.in_0011.n0 multiplexer_0.in_0011.t0 83.695
R5335 multiplexer_0.in_0011.n4 multiplexer_0.in_0011.t1 10.5295
R5336 multiplexer_0.in_0011.n4 multiplexer_0.in_0011.t2 10.5285
R5337 multiplexer_0.in_0011 multiplexer_0.in_0011.n3 4.50875
R5338 multiplexer_0.in_0011.n2 multiplexer_0.in_0011.n1 4.34635
R5339 multiplexer_0.in_0011.n1 multiplexer_0.in_0011.n0 1.5005
R5340 multiplexer_0.in_0011 multiplexer_0.in_0011.n4 0.872792
R5341 multiplexer_0.in_0011.n3 multiplexer_0.in_0011 0.177654
R5342 multiplexer_0.in_0011.n1 multiplexer_0.in_0011 0.104667
R5343 multiplexer_0.in_0011.n2 multiplexer_0.in_0011 0.0064902
R5344 multiplexer_0.in_0011.n3 multiplexer_0.in_0011.n2 0.00411538
R5345 a_n8898_n1581.t0 a_n8898_n1581.t1 21.341
R5346 a_n5142_n1581.t0 a_n5142_n1581.t1 21.167
R5347 a_n15874_1821.t0 a_n15874_1821.t1 21.2567
R5348 a_n12654_2199.t0 a_n12654_2199.t1 21.167
R5349 a_n8898_n69.t0 a_n8898_n69.t1 21.341
R5350 a_n12118_11271.t0 a_n12118_11271.t1 21.2567
R5351 multiplexer_0.in_0111.n0 multiplexer_0.in_0111.t3 228.216
R5352 multiplexer_0.in_0111.n0 multiplexer_0.in_0111.t0 83.695
R5353 multiplexer_0.in_0111.n4 multiplexer_0.in_0111.t1 10.5295
R5354 multiplexer_0.in_0111.n4 multiplexer_0.in_0111.t2 10.5285
R5355 multiplexer_0.in_0111.n2 multiplexer_0.in_0111.n1 4.34635
R5356 multiplexer_0.in_0111 multiplexer_0.in_0111.n3 4.17122
R5357 multiplexer_0.in_0111.n1 multiplexer_0.in_0111.n0 1.5005
R5358 multiplexer_0.in_0111 multiplexer_0.in_0111.n4 0.872792
R5359 multiplexer_0.in_0111.n3 multiplexer_0.in_0111 0.177654
R5360 multiplexer_0.in_0111.n1 multiplexer_0.in_0111 0.104667
R5361 multiplexer_0.in_0111.n2 multiplexer_0.in_0111 0.0064902
R5362 multiplexer_0.in_0111.n3 multiplexer_0.in_0111.n2 0.00411538
R5363 a_n15874_11649.t0 a_n15874_11649.t1 21.2567
R5364 a_n12654_12027.t0 a_n12654_12027.t1 21.167
R5365 a_n12654_8247.t0 a_n12654_8247.t1 21.167
R5366 multiplexer_0.in_1111.n0 multiplexer_0.in_1111.t3 228.216
R5367 multiplexer_0.in_1111.n0 multiplexer_0.in_1111.t0 83.695
R5368 multiplexer_0.in_1111.n4 multiplexer_0.in_1111.t1 10.5295
R5369 multiplexer_0.in_1111.n4 multiplexer_0.in_1111.t2 10.5285
R5370 multiplexer_0.in_1111.n2 multiplexer_0.in_1111.n1 4.34635
R5371 multiplexer_0.in_1111 multiplexer_0.in_1111.n3 3.28379
R5372 multiplexer_0.in_1111.n1 multiplexer_0.in_1111.n0 1.5005
R5373 multiplexer_0.in_1111 multiplexer_0.in_1111.n4 0.872792
R5374 multiplexer_0.in_1111.n3 multiplexer_0.in_1111 0.177654
R5375 multiplexer_0.in_1111.n1 multiplexer_0.in_1111 0.104667
R5376 multiplexer_0.in_1111.n2 multiplexer_0.in_1111 0.0064902
R5377 multiplexer_0.in_1111.n3 multiplexer_0.in_1111.n2 0.00411538
R5378 a_n15874_5601.t0 a_n15874_5601.t1 21.2567
R5379 multiplexer_0.trans_gate_m_25.in.t1 multiplexer_0.trans_gate_m_25.in.n0 228.216
R5380 multiplexer_0.trans_gate_m_25.in.n5 multiplexer_0.trans_gate_m_25.in.n0 1.5005
R5381 multiplexer_0.trans_gate_m_25.in.n0 multiplexer_0.trans_gate_m_25.in.t4 83.695
R5382 multiplexer_0.trans_gate_m_25.in multiplexer_0.trans_gate_m_25.in.n5 0.104667
R5383 multiplexer_0.trans_gate_m_25.in.n5 multiplexer_0.trans_gate_m_25.in.n4 4.43682
R5384 multiplexer_0.trans_gate_m_25.in.n2 multiplexer_0.trans_gate_m_25.in.n1 1.5005
R5385 multiplexer_0.trans_gate_m_25.in multiplexer_0.trans_gate_m_25.in.n2 0.104667
R5386 multiplexer_0.trans_gate_m_25.in.n4 multiplexer_0.trans_gate_m_25.in.n2 0.459875
R5387 multiplexer_0.trans_gate_m_25.in.n4 multiplexer_0.trans_gate_m_25.in 0.564042
R5388 multiplexer_0.trans_gate_m_25.in multiplexer_0.trans_gate_m_25.in.n3 1.60467
R5389 multiplexer_0.trans_gate_m_25.in.n3 multiplexer_0.trans_gate_m_25.in.t2 83.695
R5390 multiplexer_0.trans_gate_m_25.in.n3 multiplexer_0.trans_gate_m_25.in.t5 228.216
R5391 multiplexer_0.trans_gate_m_25.in.n1 multiplexer_0.trans_gate_m_25.in.t0 83.695
R5392 multiplexer_0.trans_gate_m_25.in.n1 multiplexer_0.trans_gate_m_25.in.t3 228.216
R5393 multiplexer_0.trans_gate_m_37.in.n0 multiplexer_0.trans_gate_m_37.in.t0 228.216
R5394 multiplexer_0.trans_gate_m_37.in.n0 multiplexer_0.trans_gate_m_37.in.t3 83.695
R5395 multiplexer_0.trans_gate_m_37.in.n2 multiplexer_0.trans_gate_m_37.in.n1 1.5005
R5396 multiplexer_0.trans_gate_m_37.in multiplexer_0.trans_gate_m_37.in.n2 0.104667
R5397 multiplexer_0.trans_gate_m_37.in.n5 multiplexer_0.trans_gate_m_37.in.n2 0.459875
R5398 multiplexer_0.trans_gate_m_37.in multiplexer_0.trans_gate_m_37.in.n5 0.553625
R5399 multiplexer_0.trans_gate_m_37.in multiplexer_0.trans_gate_m_37.in.n0 1.60467
R5400 multiplexer_0.trans_gate_m_37.in.n5 multiplexer_0.trans_gate_m_37.in.n4 4.43682
R5401 multiplexer_0.trans_gate_m_37.in.n4 multiplexer_0.trans_gate_m_37.in.n3 1.5005
R5402 multiplexer_0.trans_gate_m_37.in multiplexer_0.trans_gate_m_37.in.n4 0.104667
R5403 multiplexer_0.trans_gate_m_37.in.n3 multiplexer_0.trans_gate_m_37.in.t2 83.695
R5404 multiplexer_0.trans_gate_m_37.in.n3 multiplexer_0.trans_gate_m_37.in.t5 228.216
R5405 multiplexer_0.trans_gate_m_37.in.n1 multiplexer_0.trans_gate_m_37.in.t4 83.695
R5406 multiplexer_0.trans_gate_m_37.in.n1 multiplexer_0.trans_gate_m_37.in.t1 228.216
R5407 a_n12118_5223.t0 a_n12118_5223.t1 21.2567
R5408 a_n8898_5601.t0 a_n8898_5601.t1 21.167
R5409 a_n8898_n1203.t0 a_n8898_n1203.t1 21.341
R5410 a_n8898_2577.t0 a_n8898_2577.t1 21.167
R5411 a_n8362_12405.t0 a_n8362_12405.t1 21.2567
R5412 multiplexer_0.in_1000.n0 multiplexer_0.in_1000.t0 228.216
R5413 multiplexer_0.in_1000.n0 multiplexer_0.in_1000.t3 83.695
R5414 multiplexer_0.in_1000.n3 multiplexer_0.in_1000.t2 10.5739
R5415 multiplexer_0.in_1000.n3 multiplexer_0.in_1000.t1 10.5739
R5416 multiplexer_0.in_1000 multiplexer_0.in_1000.n2 3.76983
R5417 multiplexer_0.in_1000 multiplexer_0.in_1000.n3 2.20538
R5418 multiplexer_0.in_1000 multiplexer_0.in_1000.n0 1.60467
R5419 multiplexer_0.in_1000.n2 multiplexer_0.in_1000 0.471654
R5420 multiplexer_0.in_1000.n1 multiplexer_0.in_1000 0.414042
R5421 multiplexer_0.in_1000.n1 multiplexer_0.in_1000 0.0140417
R5422 multiplexer_0.in_1000.n2 multiplexer_0.in_1000.n1 0.0101154
R5423 multiplexer_0.trans_gate_m_31.in.t1 multiplexer_0.trans_gate_m_31.in.n0 228.216
R5424 multiplexer_0.trans_gate_m_31.in.n6 multiplexer_0.trans_gate_m_31.in.n0 1.5005
R5425 multiplexer_0.trans_gate_m_31.in.n0 multiplexer_0.trans_gate_m_31.in.t3 83.695
R5426 multiplexer_0.trans_gate_m_31.in multiplexer_0.trans_gate_m_31.in.n6 0.104667
R5427 multiplexer_0.trans_gate_m_31.in.n3 multiplexer_0.trans_gate_m_31.in.n4 10.4956
R5428 multiplexer_0.trans_gate_m_31.in.n3 multiplexer_0.trans_gate_m_31.in.n2 2.45249
R5429 multiplexer_0.trans_gate_m_31.in.n6 multiplexer_0.trans_gate_m_31.in.n3 2.44157
R5430 multiplexer_0.trans_gate_m_31.in.n4 multiplexer_0.trans_gate_m_31.in.n5 1.5005
R5431 multiplexer_0.trans_gate_m_31.in multiplexer_0.trans_gate_m_31.in.n4 0.104667
R5432 multiplexer_0.trans_gate_m_31.in.n5 multiplexer_0.trans_gate_m_31.in.t5 83.695
R5433 multiplexer_0.trans_gate_m_31.in.n5 multiplexer_0.trans_gate_m_31.in.t2 228.216
R5434 multiplexer_0.trans_gate_m_31.in.n2 multiplexer_0.trans_gate_m_31.in.n1 1.5005
R5435 multiplexer_0.trans_gate_m_31.in multiplexer_0.trans_gate_m_31.in.n2 0.104667
R5436 multiplexer_0.trans_gate_m_31.in.n1 multiplexer_0.trans_gate_m_31.in.t0 83.695
R5437 multiplexer_0.trans_gate_m_31.in.n1 multiplexer_0.trans_gate_m_31.in.t4 228.216
R5438 multiplexer_0.in_0001.n0 multiplexer_0.in_0001.t3 228.216
R5439 multiplexer_0.in_0001.n0 multiplexer_0.in_0001.t0 83.695
R5440 multiplexer_0.in_0001.n3 multiplexer_0.in_0001.t1 10.5295
R5441 multiplexer_0.in_0001.n3 multiplexer_0.in_0001.t2 10.5285
R5442 multiplexer_0.in_0001 multiplexer_0.in_0001.n2 4.87616
R5443 multiplexer_0.in_0001 multiplexer_0.in_0001.n0 1.60467
R5444 multiplexer_0.in_0001 multiplexer_0.in_0001.n3 0.872792
R5445 multiplexer_0.in_0001.n2 multiplexer_0.in_0001 0.471654
R5446 multiplexer_0.in_0001.n1 multiplexer_0.in_0001 0.414042
R5447 multiplexer_0.in_0001.n1 multiplexer_0.in_0001 0.0140417
R5448 multiplexer_0.in_0001.n2 multiplexer_0.in_0001.n1 0.0101154
R5449 a_n12654_n825.t0 a_n12654_n825.t1 21.341
R5450 a_n8898_n825.t0 a_n8898_n825.t1 21.34
R5451 a_n15874_9381.t0 a_n15874_9381.t1 21.2567
R5452 a_n12654_9759.t0 a_n12654_9759.t1 21.167
R5453 a_n12654_10515.t0 a_n12654_10515.t1 21.167
R5454 a_n5142_12027.t0 a_n5142_12027.t1 21.167
R5455 a_n8898_6357.t0 a_n8898_6357.t1 21.167
R5456 a_n12654_2955.t0 a_n12654_2955.t1 21.167
R5457 a_n12118_12783.t0 a_n12118_12783.t1 21.2567
R5458 a_n8898_13161.t0 a_n8898_13161.t1 21.167
R5459 a_n15874_7113.t0 a_n15874_7113.t1 21.2567
R5460 a_n12654_7491.t0 a_n12654_7491.t1 21.167
R5461 a_n15874_10137.t0 a_n15874_10137.t1 21.2567
R5462 a_n12118_3711.t0 a_n12118_3711.t1 21.2567
R5463 vtrip[3].n2 vtrip[3].t3 99.4021
R5464 vtrip[3].n0 vtrip[3].t0 23.1698
R5465 vtrip[3].n1 vtrip[3].t1 17.7681
R5466 vtrip[3].n0 vtrip[3].t2 17.7475
R5467 vtrip[3].n2 vtrip[3] 4.9564
R5468 vtrip[3].n3 vtrip[3].n2 1.7055
R5469 vtrip[3].n1 vtrip[3].n0 0.572059
R5470 vtrip[3].n3 vtrip[3].n1 0.1139
R5471 vtrip[3] vtrip[3].n3 0.0378665
R5472 a_n15874_309.t0 a_n15874_309.t1 21.2567
R5473 a_n12654_687.t0 a_n12654_687.t1 21.34
R5474 a_n12654_14295.t0 a_n12654_14295.t1 21.167
R5475 ibias.n0 ibias.t0 83.4559
R5476 ibias.n0 ibias.t1 42.9482
R5477 ibias.n1 ibias.n0 0.118921
R5478 ibias.n1 ibias 0.0613553
R5479 ibias ibias.n1 0.0605649
R5480 a_n12654_6735.t0 a_n12654_6735.t1 21.167
R5481 a_n15874_4089.t0 a_n15874_4089.t1 21.2567
R5482 a_n8898_13917.t0 a_n8898_13917.t1 21.167
R5483 level_shifter_1.in_b.n0 level_shifter_1.in_b.t1 83.7172
R5484 level_shifter_1.in_b.n0 level_shifter_1.in_b.t0 229.644
R5485 level_shifter_1.in_b level_shifter_1.in_b.n0 5.2032
R5486 level_shifter_1.in_b level_shifter_1.in_b.t2 21.9226
R5487 a_n12118_13539.t0 a_n12118_13539.t1 21.2567
R5488 a_n12654_1443.t0 a_n12654_1443.t1 21.34
R5489 a_n8898_1443.t0 a_n8898_1443.t1 21.341
R5490 a_n8362_7113.t0 a_n8362_7113.t1 21.2567
R5491 a_n12654_309.t0 a_n12654_309.t1 21.34
R5492 a_n5142_n69.t0 a_n5142_n69.t1 21.167
R5493 a_n8898_687.t0 a_n8898_687.t1 21.341
R5494 a_n8362_10893.t0 a_n8362_10893.t1 21.2567
R5495 a_n5142_11271.t0 a_n5142_11271.t1 21.167
R5496 a_n12654_n1581.t0 a_n12654_n1581.t1 21.341
R5497 a_n15874_7869.t0 a_n15874_7869.t1 21.2567
R5498 a_n8898_309.t0 a_n8898_309.t1 21.341
R5499 a_n8898_4845.t0 a_n8898_4845.t1 21.167
R5500 a_n12118_2199.t0 a_n12118_2199.t1 21.2567
R5501 a_n8898_15051.t0 a_n8898_15051.t1 21.341
R5502 a_n12118_9003.t0 a_n12118_9003.t1 21.2567
R5503 a_n12654_n1203.t0 a_n12654_n1203.t1 21.341
R5504 a_n12654_5223.t0 a_n12654_5223.t1 21.167
R5505 a_n15874_2577.t0 a_n15874_2577.t1 21.2567
R5506 a_n8898_n1959.t0 a_n8898_n1959.t1 21.341
R5507 a_n8898_12405.t0 a_n8898_12405.t1 21.167
R5508 a_n8362_7869.t0 a_n8362_7869.t1 21.2567
R5509 a_n12654_12783.t0 a_n12654_12783.t1 21.167
R5510 ovout.n0 ovout.t0 92.1108
R5511 ovout.n1 ovout.t2 83.8097
R5512 ovout ovout.n1 40.1875
R5513 ovout.n0 ovout.t1 30.088
R5514 ovout.n1 ovout.n0 1.79228
R5515 a_n8362_11649.t0 a_n8362_11649.t1 21.2567
R5516 a_n8898_8625.t0 a_n8898_8625.t1 21.167
R5517 a_n12118_5979.t0 a_n12118_5979.t1 21.2567
R5518 a_n15874_n1203.t0 a_n15874_n1203.t1 21.2567
R5519 a_n15874_13917.t0 a_n15874_13917.t1 21.2567
R5520 a_n5142_10515.t0 a_n5142_10515.t1 21.167
R5521 a_n15874_12405.t0 a_n15874_12405.t1 21.2567
C0 avss level_shifter_1.in_b 2.18706f
C1 avdd multiplexer_0.trans_gate_m_19.in 1.02912f
C2 avss multiplexer_0.in_0010 4.2278f
C3 multiplexer_0.vtrip_2 multiplexer_0.vtrip_2_b 4.73687f
C4 avss multiplexer_0.trans_gate_m_37.out 4.18674f
C5 multiplexer_0.vtrip_2_b multiplexer_0.vtrip_1_b 1.02458f
C6 ovout dvdd 1.53391f
C7 avdd multiplexer_0.trans_gate_m_18.in 1.14833f
C8 multiplexer_0.vtrip_0_b multiplexer_0.trans_gate_m_27.in 1.75429f
C9 multiplexer_0.in_1110 multiplexer_0.in_1101 1.19158f
C10 multiplexer_0.in_0110 multiplexer_0.in_0111 1.93292f
C11 avss multiplexer_0.in_1011 3.00943f
C12 vtrip[2] dvdd 3.75907f
C13 multiplexer_0.vtrip_0 multiplexer_0.trans_gate_m_23.in 1.43635f
C14 comp_hyst_0.ena_b ena 2.60102f
C15 avss multiplexer_0.in_0110 3.40355f
C16 comp_hyst_0.net1 vbg 1.36357f
C17 avss multiplexer_0.vtrip_3 5.38855f
C18 multiplexer_0.in_0000 multiplexer_0.in_0001 1.29723f
C19 ovout comp_hyst_0.net3 1.56846f
C20 multiplexer_0.trans_gate_m_37.out avdd 1.00458f
C21 avss multiplexer_0.vtrip_3_b 5.00095f
C22 vtrip[2] vtrip[3] 2.12757f
C23 avss multiplexer_0.vtrip_2 7.38242f
C24 avss multiplexer_0.vtrip_1_b 10.115201f
C25 avss multiplexer_0.vtrip_2_b 6.85919f
C26 avss multiplexer_0.in_0000 4.60989f
C27 avss multiplexer_0.trans_gate_m_21.in 2.97307f
C28 multiplexer_0.in_1011 multiplexer_0.in_1010 2.36311f
C29 avss multiplexer_0.trans_gate_m_31.out 3.01788f
C30 avss ena 8.227719f
C31 avss vin 4.26173f
C32 multiplexer_0.in_1001 multiplexer_0.in_1000 1.92146f
C33 avss multiplexer_0.trans_gate_m_33.in 4.32599f
C34 avss multiplexer_0.trans_gate_m_23.in 3.36257f
C35 avss multiplexer_0.vtrip_0 18.3412f
C36 multiplexer_0.vtrip_0_b multiplexer_0.trans_gate_m_18.in 1.67808f
C37 avss multiplexer_0.in_0111 3.37409f
C38 avdd multiplexer_0.vtrip_3 5.64672f
C39 multiplexer_0.vtrip_3_b avdd 3.56297f
C40 avss vtrip[1] 1.94321f
C41 multiplexer_0.vtrip_2 avdd 11.521f
C42 avss multiplexer_0.in_0001 3.89824f
C43 multiplexer_0.vtrip_1_b avdd 10.187099f
C44 avss multiplexer_0.in_0100 3.71413f
C45 multiplexer_0.vtrip_2_b avdd 6.36948f
C46 multiplexer_0.trans_gate_m_21.in avdd 1.04208f
C47 multiplexer_0.in_1101 multiplexer_0.in_1100 1.47135f
C48 multiplexer_0.trans_gate_m_31.out avdd 1.14658f
C49 avdd vin 1.31175f
C50 multiplexer_0.trans_gate_m_33.in avdd 1.31623f
C51 multiplexer_0.trans_gate_m_32.in multiplexer_0.vtrip_2 1.03862f
C52 multiplexer_0.vtrip_0 avdd 22.856901f
C53 multiplexer_0.trans_gate_m_23.in avdd 1.15181f
C54 multiplexer_0.in_0011 multiplexer_0.in_0010 2.38759f
C55 ena dvdd 5.53155f
C56 vin dvdd 1.15918f
C57 multiplexer_0.vtrip_1_b multiplexer_0.vtrip_1 7.7058f
C58 level_shifter_2.in_b vtrip[2] 2.32089f
C59 vbg vin 2.9135f
C60 comp_hyst_0.ena_b dvdd 2.6983f
C61 vtrip[1] dvdd 3.94954f
C62 multiplexer_0.vtrip_2 multiplexer_0.trans_gate_m_28.in 1.01863f
C63 avss avdd 1.62977p
C64 avss multiplexer_0.in_1111 3.34253f
C65 avss multiplexer_0.in_1010 2.8365f
C66 avss level_shifter_0.in_b 1.92248f
C67 multiplexer_0.in_0110 multiplexer_0.in_0011 1.4217f
C68 comp_hyst_0.net5 comp_hyst_0.net1 2.80231f
C69 multiplexer_0.vtrip_0 multiplexer_0.trans_gate_m_31.in 1.42693f
C70 avss multiplexer_0.in_1110 2.8304f
C71 avss multiplexer_0.trans_gate_m_32.in 2.96668f
C72 avss multiplexer_0.vtrip_1 11.345901f
C73 multiplexer_0.vtrip_0 multiplexer_0.trans_gate_m_27.in 1.45603f
C74 avss vtrip[3] 2.52607f
C75 avss multiplexer_0.trans_gate_m_29.in 3.01849f
C76 comp_hyst_0.net2 comp_hyst_0.net4 1.09495f
C77 multiplexer_0.vtrip_0_b multiplexer_0.trans_gate_m_23.in 1.56933f
C78 multiplexer_0.vtrip_0 multiplexer_0.vtrip_0_b 8.32478f
C79 vtrip[0] vtrip[1] 3.22357f
C80 avss multiplexer_0.trans_gate_m_28.in 2.85568f
C81 avss multiplexer_0.trans_gate_m_31.in 3.40808f
C82 avss multiplexer_0.trans_gate_m_25.in 2.91806f
C83 multiplexer_0.in_1111 multiplexer_0.in_1110 1.60188f
C84 avss vtrip[0] 1.54546f
C85 multiplexer_0.trans_gate_m_32.in avdd 1.02713f
C86 multiplexer_0.vtrip_1 avdd 17.3142f
C87 multiplexer_0.in_0110 multiplexer_0.in_0101 1.83216f
C88 avss multiplexer_0.trans_gate_m_27.in 3.34445f
C89 avss multiplexer_0.vtrip_0_b 15.788701f
C90 multiplexer_0.trans_gate_m_29.in avdd 1.03758f
C91 avss multiplexer_0.in_0011 3.46624f
C92 vtrip[3] dvdd 2.30283f
C93 avss level_shifter_3.in_b 2.22418f
C94 comp_hyst_0.net4 dvdd 30.420599f
C95 ibias dvdd 4.8744f
C96 avdd multiplexer_0.trans_gate_m_28.in 1.01616f
C97 avss multiplexer_0.in_1001 2.85342f
C98 multiplexer_0.trans_gate_m_31.in avdd 1.15303f
C99 comp_hyst_0.net5 ena 1.53335f
C100 multiplexer_0.in_0111 multiplexer_0.in_1000 1.1086f
C101 vbg comp_hyst_0.net4 1.89072f
C102 comp_hyst_0.net3 dvdd 45.820198f
C103 avdd multiplexer_0.trans_gate_m_25.in 1.02269f
C104 avss multiplexer_0.in_1100 2.55289f
C105 vbg comp_hyst_0.net3 1.08435f
C106 multiplexer_0.vtrip_0 multiplexer_0.trans_gate_m_18.in 1.42669f
C107 comp_hyst_0.ena_b comp_hyst_0.net5 2.09269f
C108 level_shifter_0.in_b vtrip[0] 2.23942f
C109 vtrip[0] dvdd 5.49537f
C110 avss level_shifter_2.in_b 2.18802f
C111 avdd multiplexer_0.trans_gate_m_27.in 1.12621f
C112 avss multiplexer_0.in_1000 3.15058f
C113 multiplexer_0.vtrip_0_b avdd 16.2951f
C114 multiplexer_0.trans_gate_m_37.out multiplexer_0.vtrip_3 1.58056f
C115 avss multiplexer_0.trans_gate_m_37.in 3.15158f
C116 comp_hyst_0.net1 vin 1.08144f
C117 multiplexer_0.in_0100 multiplexer_0.in_0101 1.4247f
C118 comp_hyst_0.net3 comp_hyst_0.net4 17.705801f
C119 avss multiplexer_0.trans_gate_m_19.in 3.04297f
C120 avss multiplexer_0.in_0101 3.35968f
C121 multiplexer_0.in_1010 multiplexer_0.in_1001 1.33401f
C122 vtrip[1] vtrip[2] 2.74924f
C123 comp_hyst_0.net2 ovout 1.14594f
C124 avss multiplexer_0.in_1101 3.55535f
C125 multiplexer_0.vtrip_0_b multiplexer_0.vtrip_1 1.91482f
C126 avss multiplexer_0.trans_gate_m_18.in 3.39154f
C127 avss vtrip[2] 2.04916f
C128 level_shifter_1.in_b vtrip[1] 2.27942f
C129 multiplexer_0.in_1010 multiplexer_0.in_1000 1.21062f
C130 level_shifter_3.in_b vtrip[3] 2.36959f
C131 avdd multiplexer_0.trans_gate_m_37.in 1.01954f
C132 multiplexer_0.vtrip_3_b multiplexer_0.vtrip_3 3.3491f
C133 multiplexer_0.trans_gate_m_31.in multiplexer_0.vtrip_0_b 1.67382f
C134 vbg dvss 11.814878f
C135 ovout dvss 4.14261f
C136 ibias dvss 9.874781f
C137 ena dvss 20.711246f
C138 vtrip[3] dvss 7.803799f
C139 vtrip[2] dvss 9.231338f
C140 vtrip[1] dvss 9.753779f
C141 vtrip[0] dvss 10.507146f
C142 avss dvss 0.406581p
C143 dvdd dvss 1.216993p
C144 avdd dvss 2.03821p
C145 m1_21598_448# dvss 4.41071f $ **FLOATING
C146 comp_hyst_0.net1 dvss 4.679739f
C147 comp_hyst_0.net5 dvss 25.12681f
C148 comp_hyst_0.net2 dvss 7.539189f
C149 comp_hyst_0.ena_b dvss 10.262756f
C150 level_shifter_3.in_b dvss 3.88048f
C151 level_shifter_2.in_b dvss 3.70586f
C152 level_shifter_1.in_b dvss 3.73365f
C153 level_shifter_0.in_b dvss 2.63882f
C154 multiplexer_0.vtrip_3_b dvss 7.874678f
C155 vin dvss 19.093369f
C156 multiplexer_0.vtrip_3 dvss 8.414051f
C157 comp_hyst_0.net3 dvss 21.120062f
C158 comp_hyst_0.net4 dvss 13.7459f
C159 multiplexer_0.vtrip_2_b dvss 7.151894f
C160 multiplexer_0.vtrip_2 dvss 7.901592f
C161 multiplexer_0.vtrip_1_b dvss 5.897985f
C162 multiplexer_0.vtrip_1 dvss 11.941719f
C163 multiplexer_0.vtrip_0_b dvss 9.68784f
C164 multiplexer_0.vtrip_0 dvss 15.1825f
C165 multiplexer_0.in_1111 dvss 1.823567f
C166 multiplexer_0.in_1110 dvss 2.124716f
C167 multiplexer_0.in_1101 dvss 1.810742f
C168 multiplexer_0.in_1100 dvss 1.583226f
C169 multiplexer_0.in_1011 dvss 2.71753f
C170 multiplexer_0.in_1010 dvss 2.890666f
C171 multiplexer_0.in_1001 dvss 1.689299f
C172 multiplexer_0.in_1000 dvss 2.181204f
C173 multiplexer_0.in_0111 dvss 1.826988f
C174 multiplexer_0.in_0110 dvss 1.901118f
C175 multiplexer_0.in_0101 dvss 2.265734f
C176 multiplexer_0.in_0100 dvss 2.550706f
C177 multiplexer_0.in_0011 dvss 2.577745f
C178 multiplexer_0.in_0010 dvss 3.263069f
C179 multiplexer_0.in_0001 dvss 1.934929f
C180 multiplexer_0.in_0000 dvss 2.276361f
C181 level_shifter_1.in_b.n0 dvss 1.15334f
C182 level_shifter_1.in_b.t2 dvss 1.11724f
C183 vtrip[3].n0 dvss 1.65578f
C184 vtrip[3].n1 dvss 2.1534f
C185 multiplexer_0.in_0001.n3 dvss 1.76738f
C186 multiplexer_0.trans_gate_m_31.in.n3 dvss 1.61117f
C187 multiplexer_0.in_1000.n3 dvss 1.48678f
C188 multiplexer_0.in_1111.n4 dvss 1.52623f
C189 multiplexer_0.in_0111.n4 dvss 1.31558f
C190 multiplexer_0.in_0011.n4 dvss 2.24729f
C191 multiplexer_0.in_1110.n4 dvss 1.30461f
C192 multiplexer_0.trans_gate_m_18.in.n3 dvss 1.61117f
C193 level_shifter_2.in_b.n0 dvss 1.15334f
C194 level_shifter_2.in_b.t2 dvss 1.11724f
C195 vtrip[2].t2 dvss 1.21331f
C196 vtrip[2].n0 dvss 2.06705f
C197 vtrip[2].n1 dvss 2.68828f
C198 vtrip[2].n2 dvss 1.29487f
C199 comp_hyst_0.ena_b.n7 dvss 1.16035f
C200 comp_hyst_0.ena_b.t5 dvss 1.74723f
C201 multiplexer_0.in_1010.n4 dvss 2.19323f
C202 multiplexer_0.trans_gate_m_33.in.n2 dvss 1.31038f
C203 multiplexer_0.trans_gate_m_33.in.n3 dvss 1.49028f
C204 multiplexer_0.vtrip_3_b.n1 dvss 1.14654f
C205 multiplexer_0.vtrip_3_b.n2 dvss 1.53645f
C206 a_n5142_n1959.t1 dvss 2.3994f
C207 ena.n5 dvss 1.0283f
C208 ena.n10 dvss 5.0478f
C209 ena.n11 dvss 2.97276f
C210 multiplexer_0.trans_gate_m_27.in.n3 dvss 1.56379f
C211 multiplexer_0.in_0101.n3 dvss 1.5916f
C212 multiplexer_0.in_0100.n3 dvss 1.6941f
C213 vbg.n0 dvss 1.25899f
C214 multiplexer_0.vtrip_2_b.n3 dvss 1.02684f
C215 multiplexer_0.vtrip_2_b.n5 dvss 1.30183f
C216 multiplexer_0.vtrip_2_b.n6 dvss 2.45453f
C217 multiplexer_0.vtrip_2_b.n7 dvss 1.57666f
C218 multiplexer_0.trans_gate_m_23.in.n3 dvss 1.61117f
C219 multiplexer_0.in_1001.n2 dvss 1.3732f
C220 vin.n3 dvss 1.76099f
C221 multiplexer_0.in_0000.n3 dvss 2.01807f
C222 multiplexer_0.vtrip_0_b.n2 dvss 1.40158f
C223 multiplexer_0.vtrip_0_b.n4 dvss 1.40616f
C224 multiplexer_0.vtrip_0_b.n7 dvss 1.40158f
C225 multiplexer_0.vtrip_0_b.n9 dvss 1.40616f
C226 multiplexer_0.vtrip_0_b.n11 dvss 1.27162f
C227 multiplexer_0.vtrip_0_b.n12 dvss 1.40158f
C228 multiplexer_0.vtrip_0_b.n14 dvss 1.40616f
C229 multiplexer_0.vtrip_0_b.n16 dvss 1.9554f
C230 multiplexer_0.vtrip_0_b.n17 dvss 1.40158f
C231 multiplexer_0.vtrip_0_b.n19 dvss 1.40616f
C232 multiplexer_0.vtrip_0_b.n21 dvss 1.67384f
C233 multiplexer_0.vtrip_0_b.n23 dvss 2.6433f
C234 multiplexer_0.vtrip_0_b.n24 dvss 2.78781f
C235 multiplexer_0.in_0010.n4 dvss 2.44947f
C236 comp_hyst_0.net1.n2 dvss 1.16757f
C237 comp_hyst_0.net5.t5 dvss 1.46711f
C238 vtrip[1].t0 dvss 1.03496f
C239 vtrip[1].n0 dvss 1.76321f
C240 vtrip[1].n1 dvss 2.29313f
C241 vtrip[1].n2 dvss 1.48872f
C242 multiplexer_0.in_1011.n3 dvss 2.20748f
C243 multiplexer_0.vtrip_0.n0 dvss 1.36646f
C244 multiplexer_0.vtrip_0.n1 dvss 1.25223f
C245 multiplexer_0.vtrip_0.n2 dvss 1.99048f
C246 multiplexer_0.vtrip_0.n3 dvss 1.72856f
C247 multiplexer_0.vtrip_0.n5 dvss 1.73422f
C248 multiplexer_0.vtrip_0.n7 dvss 2.02902f
C249 multiplexer_0.vtrip_0.n8 dvss 1.72856f
C250 multiplexer_0.vtrip_0.n10 dvss 1.73422f
C251 multiplexer_0.vtrip_0.n12 dvss 1.00107f
C252 multiplexer_0.vtrip_0.n13 dvss 1.72856f
C253 multiplexer_0.vtrip_0.n15 dvss 1.73422f
C254 multiplexer_0.vtrip_0.t10 dvss 1.01084f
C255 multiplexer_0.vtrip_0.n18 dvss 1.01955f
C256 multiplexer_0.vtrip_0.t3 dvss 1.0194f
C257 multiplexer_0.vtrip_0.n20 dvss 1.13693f
C258 multiplexer_0.vtrip_0.n23 dvss 1.20822f
C259 multiplexer_0.vtrip_0.n24 dvss 2.93945f
C260 avdd.n1 dvss 5.39489f
C261 avdd.n3 dvss 5.39489f
C262 avdd.t5 dvss 7.22231f
C263 avdd.n9 dvss 2.06399f
C264 avdd.n10 dvss 1.72384f
C265 avdd.n12 dvss 5.39489f
C266 avdd.n14 dvss 5.39489f
C267 avdd.t16 dvss 7.22231f
C268 avdd.n20 dvss 2.06399f
C269 avdd.n21 dvss 1.72384f
C270 avdd.n23 dvss 5.39489f
C271 avdd.n25 dvss 5.39489f
C272 avdd.t7 dvss 7.22231f
C273 avdd.n31 dvss 2.06399f
C274 avdd.n32 dvss 1.72384f
C275 avdd.n34 dvss 5.39489f
C276 avdd.n36 dvss 5.39489f
C277 avdd.t35 dvss 7.22231f
C278 avdd.n42 dvss 2.06399f
C279 avdd.n43 dvss 1.72384f
C280 avdd.n45 dvss 5.39489f
C281 avdd.n47 dvss 5.39489f
C282 avdd.t33 dvss 7.22231f
C283 avdd.n53 dvss 2.06399f
C284 avdd.n54 dvss 1.72384f
C285 avdd.n56 dvss 5.39489f
C286 avdd.n58 dvss 5.39489f
C287 avdd.t10 dvss 7.22231f
C288 avdd.n64 dvss 2.06399f
C289 avdd.n65 dvss 1.72384f
C290 avdd.n67 dvss 5.39489f
C291 avdd.n69 dvss 5.39489f
C292 avdd.t15 dvss 7.22231f
C293 avdd.n75 dvss 2.06399f
C294 avdd.n76 dvss 1.72384f
C295 avdd.n78 dvss 5.39489f
C296 avdd.n80 dvss 5.39489f
C297 avdd.t0 dvss 7.22231f
C298 avdd.n86 dvss 2.06399f
C299 avdd.n87 dvss 1.72384f
C300 avdd.n89 dvss 5.39489f
C301 avdd.n91 dvss 5.39489f
C302 avdd.t26 dvss 7.22231f
C303 avdd.n97 dvss 2.06399f
C304 avdd.n98 dvss 1.72384f
C305 avdd.n100 dvss 5.39489f
C306 avdd.n102 dvss 5.39489f
C307 avdd.t9 dvss 7.22231f
C308 avdd.n108 dvss 2.06399f
C309 avdd.n109 dvss 1.72384f
C310 avdd.n111 dvss 5.39489f
C311 avdd.n113 dvss 5.39489f
C312 avdd.t12 dvss 7.22231f
C313 avdd.n119 dvss 2.06399f
C314 avdd.n120 dvss 1.72384f
C315 avdd.n122 dvss 5.39489f
C316 avdd.n124 dvss 5.39489f
C317 avdd.t6 dvss 7.22231f
C318 avdd.n130 dvss 2.06399f
C319 avdd.n131 dvss 1.72384f
C320 avdd.n133 dvss 5.39489f
C321 avdd.n135 dvss 5.39489f
C322 avdd.t4 dvss 7.22231f
C323 avdd.n141 dvss 2.06399f
C324 avdd.n142 dvss 1.72384f
C325 avdd.n144 dvss 5.39489f
C326 avdd.n146 dvss 5.39489f
C327 avdd.t34 dvss 7.22231f
C328 avdd.n152 dvss 2.06399f
C329 avdd.n153 dvss 1.72384f
C330 avdd.n155 dvss 5.39489f
C331 avdd.n157 dvss 5.39489f
C332 avdd.t17 dvss 7.22231f
C333 avdd.n163 dvss 2.06399f
C334 avdd.n164 dvss 1.72384f
C335 avdd.n166 dvss 5.39489f
C336 avdd.n168 dvss 5.39489f
C337 avdd.t8 dvss 7.22231f
C338 avdd.n174 dvss 2.06399f
C339 avdd.n175 dvss 1.72384f
C340 avdd.n177 dvss 5.39489f
C341 avdd.n179 dvss 5.39489f
C342 avdd.t38 dvss 7.22231f
C343 avdd.n185 dvss 2.06399f
C344 avdd.n186 dvss 1.72384f
C345 avdd.n188 dvss 5.39489f
C346 avdd.n190 dvss 5.39489f
C347 avdd.t22 dvss 7.22231f
C348 avdd.n196 dvss 2.06399f
C349 avdd.n197 dvss 1.72384f
C350 avdd.n199 dvss 5.39489f
C351 avdd.n201 dvss 5.39489f
C352 avdd.t40 dvss 7.22231f
C353 avdd.n207 dvss 2.06399f
C354 avdd.n208 dvss 1.72384f
C355 avdd.n210 dvss 5.39489f
C356 avdd.n212 dvss 5.39489f
C357 avdd.t23 dvss 7.22231f
C358 avdd.n218 dvss 2.06399f
C359 avdd.n219 dvss 1.72384f
C360 avdd.n221 dvss 5.39489f
C361 avdd.n223 dvss 5.39489f
C362 avdd.t36 dvss 7.22231f
C363 avdd.n229 dvss 2.06399f
C364 avdd.n230 dvss 1.72384f
C365 avdd.n232 dvss 5.39489f
C366 avdd.n234 dvss 5.39489f
C367 avdd.t20 dvss 7.22231f
C368 avdd.n240 dvss 2.06399f
C369 avdd.n241 dvss 1.72384f
C370 avdd.n243 dvss 5.39489f
C371 avdd.n245 dvss 5.39489f
C372 avdd.t37 dvss 7.22231f
C373 avdd.n251 dvss 2.06399f
C374 avdd.n252 dvss 1.72384f
C375 avdd.n254 dvss 5.39489f
C376 avdd.n256 dvss 5.39489f
C377 avdd.t21 dvss 7.22231f
C378 avdd.n262 dvss 2.06399f
C379 avdd.n263 dvss 1.72384f
C380 avdd.n265 dvss 5.39489f
C381 avdd.n267 dvss 5.39489f
C382 avdd.t3 dvss 7.22231f
C383 avdd.n273 dvss 2.06399f
C384 avdd.n274 dvss 3.44767f
C385 avdd.n276 dvss 5.39489f
C386 avdd.n278 dvss 5.39489f
C387 avdd.t31 dvss 7.22231f
C388 avdd.n284 dvss 2.06399f
C389 avdd.n285 dvss 1.72384f
C390 avdd.n287 dvss 5.39489f
C391 avdd.n289 dvss 5.39489f
C392 avdd.t11 dvss 7.22231f
C393 avdd.n295 dvss 2.06399f
C394 avdd.n296 dvss 3.44767f
C395 avdd.n298 dvss 5.39489f
C396 avdd.n300 dvss 5.39489f
C397 avdd.t30 dvss 7.22231f
C398 avdd.n306 dvss 2.06399f
C399 avdd.n307 dvss 1.72384f
C400 avdd.n308 dvss 2.802f
C401 avdd.n313 dvss 8.426219f
C402 avdd.n315 dvss 8.426219f
C403 avdd.n325 dvss 9.74957f
C404 avdd.t24 dvss 11.948999f
C405 avdd.n328 dvss 1.93421f
C406 avdd.n329 dvss 2.93397f
C407 avdd.n330 dvss 2.80158f
C408 avdd.n331 dvss 2.802f
C409 avdd.n336 dvss 8.426219f
C410 avdd.n338 dvss 8.426219f
C411 avdd.n348 dvss 9.74957f
C412 avdd.t1 dvss 11.948999f
C413 avdd.n351 dvss 1.93421f
C414 avdd.n352 dvss 2.93397f
C415 avdd.n353 dvss 2.80158f
C416 avdd.n354 dvss 8.42617f
C417 avdd.n355 dvss 2.802f
C418 avdd.n360 dvss 8.426219f
C419 avdd.n362 dvss 8.426219f
C420 avdd.n372 dvss 9.74957f
C421 avdd.t18 dvss 11.948999f
C422 avdd.n375 dvss 1.93421f
C423 avdd.n376 dvss 2.93397f
C424 avdd.n377 dvss 2.80158f
C425 avdd.n378 dvss 8.02315f
C426 avdd.n379 dvss 2.802f
C427 avdd.n384 dvss 8.426219f
C428 avdd.n386 dvss 8.426219f
C429 avdd.n396 dvss 9.74957f
C430 avdd.t13 dvss 11.948999f
C431 avdd.n399 dvss 1.93421f
C432 avdd.n400 dvss 2.93397f
C433 avdd.n401 dvss 2.80158f
C434 avdd.n402 dvss 24.6949f
C435 avdd.n403 dvss 0.105131p
C436 avdd.n404 dvss 46.7712f
C437 avdd.n405 dvss 46.327503f
C438 avdd.n406 dvss 63.9731f
C439 avdd.n407 dvss 13.3624f
C440 avdd.n408 dvss 0.20923p
C441 multiplexer_0.trans_gate_m_37.out.n4 dvss 1.45563f
C442 multiplexer_0.trans_gate_m_37.out.n5 dvss 1.27991f
C443 vtrip[0].n0 dvss 1.45751f
C444 vtrip[0].n1 dvss 1.89554f
C445 vtrip[0].n2 dvss 1.6207f
C446 multiplexer_0.in_1101.n3 dvss 1.7658f
C447 multiplexer_0.in_1100.n3 dvss 1.37623f
C448 multiplexer_0.vtrip_2.n0 dvss 1.52182f
C449 multiplexer_0.vtrip_2.n1 dvss 1.3946f
C450 multiplexer_0.vtrip_2.t6 dvss 1.09443f
C451 multiplexer_0.vtrip_2.t7 dvss 1.09421f
C452 multiplexer_0.vtrip_2.n2 dvss 1.82632f
C453 multiplexer_0.vtrip_2.t4 dvss 1.1353f
C454 multiplexer_0.vtrip_2.n3 dvss 1.82127f
C455 multiplexer_0.vtrip_2.n4 dvss 1.93139f
C456 multiplexer_0.vtrip_2.t5 dvss 1.00389f
C457 multiplexer_0.vtrip_2.t3 dvss 1.04296f
C458 multiplexer_0.vtrip_2.n5 dvss 1.04904f
C459 multiplexer_0.vtrip_2.n6 dvss 3.38267f
C460 multiplexer_0.in_0110.n4 dvss 1.28133f
C461 multiplexer_0.vtrip_3.n0 dvss 1.35303f
C462 multiplexer_0.vtrip_3.n1 dvss 1.23992f
C463 multiplexer_0.vtrip_3.t5 dvss 1.00938f
C464 multiplexer_0.vtrip_3.n3 dvss 1.53947f
C465 level_shifter_3.in_b.n0 dvss 1.17897f
C466 level_shifter_3.in_b.t2 dvss 1.14207f
C467 comp_hyst_0.net3.n0 dvss 1.22259f
C468 comp_hyst_0.net3.n1 dvss 2.52721f
C469 comp_hyst_0.net3.n2 dvss 1.52394f
C470 comp_hyst_0.net3.n3 dvss 2.40127f
C471 comp_hyst_0.net3.t10 dvss 3.5614f
C472 comp_hyst_0.net3.n4 dvss 1.52394f
C473 comp_hyst_0.net3.t6 dvss 3.51069f
C474 comp_hyst_0.net3.n6 dvss 2.40127f
C475 comp_hyst_0.net3.t9 dvss 6.06936f
C476 comp_hyst_0.net3.n7 dvss 2.63343f
C477 comp_hyst_0.net3.n8 dvss 2.633f
C478 comp_hyst_0.net3.n11 dvss 1.52394f
C479 comp_hyst_0.net3.n12 dvss 2.40127f
C480 comp_hyst_0.net3.t13 dvss 3.5614f
C481 comp_hyst_0.net3.n13 dvss 1.52394f
C482 comp_hyst_0.net3.t4 dvss 3.51069f
C483 comp_hyst_0.net3.n15 dvss 2.40127f
C484 comp_hyst_0.net3.t11 dvss 6.06936f
C485 comp_hyst_0.net3.n16 dvss 2.633f
C486 comp_hyst_0.net3.n17 dvss 2.633f
C487 comp_hyst_0.net3.n20 dvss 2.28622f
C488 dvdd.n50 dvss 2.59665f
C489 dvdd.n51 dvss 1.29818f
C490 dvdd.n52 dvss 1.40778f
C491 dvdd.n55 dvss 2.85795f
C492 dvdd.n56 dvss 2.85795f
C493 dvdd.n70 dvss 1.6282f
C494 dvdd.n97 dvss 1.6282f
C495 dvdd.n134 dvss 1.43542f
C496 dvdd.n135 dvss 1.43542f
C497 dvdd.t6 dvss 2.28264f
C498 dvdd.n421 dvss 1.52361f
C499 dvdd.n424 dvss 12.7602f
C500 dvdd.n425 dvss 1.35293f
C501 dvdd.n478 dvss 1.49529f
C502 dvdd.n479 dvss 1.27502f
C503 dvdd.n620 dvss 1.40467f
C504 dvdd.t16 dvss 2.85795f
C505 dvdd.n652 dvss 1.40467f
C506 dvdd.t18 dvss 2.85795f
C507 dvdd.t13 dvss 2.85795f
C508 dvdd.n662 dvss 3.31573f
C509 dvdd.n663 dvss 14.948f
C510 dvdd.n664 dvss 5.33263f
C511 dvdd.n665 dvss 2.76314f
C512 dvdd.n667 dvss 1.10126f
C513 comp_hyst_0.net4.t13 dvss 3.2071f
C514 comp_hyst_0.net4.n1 dvss 1.28102f
C515 comp_hyst_0.net4.n5 dvss 1.69638f
C516 comp_hyst_0.net4.t3 dvss 2.25721f
C517 comp_hyst_0.net4.n6 dvss 1.53524f
C518 comp_hyst_0.net4.n9 dvss 1.69638f
C519 comp_hyst_0.net4.n11 dvss 1.53568f
C520 comp_hyst_0.net4.t1 dvss 2.25707f
C521 comp_hyst_0.net4.n12 dvss 1.32518f
C522 comp_hyst_0.net4.n13 dvss 1.51759f
C523 comp_hyst_0.net4.t11 dvss 3.20661f
C524 comp_hyst_0.net4.n14 dvss 1.80073f
C525 comp_hyst_0.net4.n15 dvss 1.47286f
C526 comp_hyst_0.net4.n16 dvss 1.47256f
C527 comp_hyst_0.net4.n17 dvss 1.69922f
C528 comp_hyst_0.net4.n21 dvss 1.54046f
C529 comp_hyst_0.net4.n22 dvss 3.58022f
C530 comp_hyst_0.net4.n24 dvss 4.70385f
C531 comp_hyst_0.net4.t12 dvss 3.56478f
C532 multiplexer_0.vtrip_1_b.n2 dvss 1.40035f
C533 multiplexer_0.vtrip_1_b.n3 dvss 1.64459f
C534 multiplexer_0.vtrip_1_b.n4 dvss 1.40035f
C535 multiplexer_0.vtrip_1_b.n5 dvss 1.06739f
C536 multiplexer_0.vtrip_1_b.n6 dvss 1.40035f
C537 multiplexer_0.vtrip_1_b.n7 dvss 1.98904f
C538 multiplexer_0.vtrip_1_b.n8 dvss 1.40035f
C539 multiplexer_0.vtrip_1_b.n9 dvss 1.31534f
C540 multiplexer_0.vtrip_1_b.n11 dvss 2.66714f
C541 multiplexer_0.vtrip_1_b.n12 dvss 3.13377f
C542 avss.n0 dvss 1.30263f
C543 avss.n1 dvss 1.88827f
C544 avss.n2 dvss 1.88849f
C545 avss.n4 dvss 1.38053f
C546 avss.n5 dvss 1.9273f
C547 avss.n6 dvss 2.12999f
C548 avss.n7 dvss 2.12999f
C549 avss.n8 dvss 2.12999f
C550 avss.n9 dvss 2.12999f
C551 avss.n10 dvss 2.12999f
C552 avss.n11 dvss 2.12999f
C553 avss.n12 dvss 2.12999f
C554 avss.n13 dvss 2.12999f
C555 avss.n14 dvss 2.12999f
C556 avss.n15 dvss 2.12999f
C557 avss.n16 dvss 2.12999f
C558 avss.n17 dvss 2.12999f
C559 avss.n18 dvss 2.12999f
C560 avss.n19 dvss 2.12999f
C561 avss.n20 dvss 2.12999f
C562 avss.n21 dvss 2.12999f
C563 avss.n22 dvss 2.12999f
C564 avss.n23 dvss 2.12999f
C565 avss.n24 dvss 2.12999f
C566 avss.n25 dvss 2.12999f
C567 avss.n26 dvss 2.12999f
C568 avss.n27 dvss 2.12999f
C569 avss.n28 dvss 2.12999f
C570 avss.n29 dvss 2.12999f
C571 avss.n30 dvss 2.12999f
C572 avss.n31 dvss 2.12999f
C573 avss.n32 dvss 2.12999f
C574 avss.n33 dvss 2.12999f
C575 avss.n34 dvss 2.12999f
C576 avss.n35 dvss 2.12999f
C577 avss.n36 dvss 2.12999f
C578 avss.n37 dvss 2.12999f
C579 avss.n38 dvss 2.12999f
C580 avss.n39 dvss 2.12999f
C581 avss.n40 dvss 2.12999f
C582 avss.n41 dvss 2.12999f
C583 avss.n42 dvss 2.12999f
C584 avss.n43 dvss 2.12999f
C585 avss.n44 dvss 2.12999f
C586 avss.n45 dvss 2.12999f
C587 avss.n46 dvss 2.12999f
C588 avss.n47 dvss 2.12999f
C589 avss.n48 dvss 2.12999f
C590 avss.n49 dvss 2.12999f
C591 avss.n50 dvss 2.12999f
C592 avss.n51 dvss 2.10879f
C593 avss.n52 dvss 1.80989f
C594 avss.n53 dvss 1.88827f
C595 avss.n54 dvss 1.88849f
C596 avss.n55 dvss 1.88827f
C597 avss.n56 dvss 1.88849f
C598 avss.n57 dvss 1.80931f
C599 avss.n58 dvss 2.10843f
C600 avss.n59 dvss 2.12999f
C601 avss.n60 dvss 2.12999f
C602 avss.n61 dvss 2.12999f
C603 avss.n62 dvss 2.12999f
C604 avss.n63 dvss 2.12999f
C605 avss.n64 dvss 2.12999f
C606 avss.n65 dvss 2.12999f
C607 avss.n66 dvss 2.12999f
C608 avss.n67 dvss 2.12999f
C609 avss.n68 dvss 2.12999f
C610 avss.n69 dvss 2.12999f
C611 avss.n70 dvss 2.12999f
C612 avss.n71 dvss 2.12999f
C613 avss.n72 dvss 2.12999f
C614 avss.n73 dvss 2.12999f
C615 avss.n74 dvss 2.12999f
C616 avss.n75 dvss 2.12999f
C617 avss.n76 dvss 2.12999f
C618 avss.n77 dvss 2.12999f
C619 avss.n78 dvss 2.12999f
C620 avss.n79 dvss 2.12999f
C621 avss.n80 dvss 2.12999f
C622 avss.n81 dvss 2.12999f
C623 avss.n82 dvss 2.12999f
C624 avss.n83 dvss 2.12999f
C625 avss.n84 dvss 2.12999f
C626 avss.n85 dvss 2.12999f
C627 avss.n86 dvss 2.12999f
C628 avss.n87 dvss 2.12999f
C629 avss.n88 dvss 2.12999f
C630 avss.n89 dvss 2.12999f
C631 avss.n90 dvss 2.12999f
C632 avss.n91 dvss 2.12999f
C633 avss.n92 dvss 2.12999f
C634 avss.n93 dvss 2.12999f
C635 avss.n94 dvss 2.12999f
C636 avss.n95 dvss 2.12999f
C637 avss.n96 dvss 2.12999f
C638 avss.n97 dvss 2.12999f
C639 avss.n98 dvss 2.12999f
C640 avss.n99 dvss 2.12999f
C641 avss.n100 dvss 2.12999f
C642 avss.n101 dvss 2.12999f
C643 avss.n102 dvss 2.12999f
C644 avss.n103 dvss 2.12999f
C645 avss.n104 dvss 1.9273f
C646 avss.n105 dvss 1.37998f
C647 avss.n107 dvss 1.88827f
C648 avss.n108 dvss 1.88849f
C649 avss.n109 dvss 1.30278f
C650 avss.n110 dvss 37.6986f
C651 avss.n111 dvss 9.978429f
C652 avss.n112 dvss 6.26811f
C653 avss.n113 dvss 2.40542f
C654 avss.n114 dvss 58.557697f
C655 avss.t0 dvss 37.5956f
C656 avss.t5 dvss 86.8916f
C657 avss.n119 dvss 15.6291f
C658 avss.t13 dvss 86.8916f
C659 avss.t14 dvss 47.4543f
C660 avss.n120 dvss 21.4327f
C661 avss.n121 dvss 15.521199f
C662 avss.n128 dvss 1.12574f
C663 avss.t31 dvss 5.01586f
C664 avss.n137 dvss 6.15944f
C665 avss.n161 dvss 18.7238f
C666 avss.n162 dvss 9.93295f
C667 avss.t41 dvss 3.84754f
C668 avss.n167 dvss 2.75401f
C669 avss.n168 dvss 3.27009f
C670 avss.t26 dvss 2.8988f
C671 avss.n206 dvss 2.62332f
C672 avss.n213 dvss 2.61079f
C673 avss.n214 dvss 3.15651f
C674 avss.n215 dvss 1.06406f
C675 avss.t60 dvss 7.624569f
C676 avss.n224 dvss 6.86705f
C677 avss.n225 dvss 3.43526f
C678 avss.n235 dvss 1.94342f
C679 avss.n239 dvss 1.94342f
C680 avss.n249 dvss 1.33105f
C681 avss.n253 dvss 1.80693f
C682 avss.n264 dvss 4.1063f
C683 avss.t158 dvss 5.7008f
C684 avss.n272 dvss 1.37613f
C685 avss.t215 dvss 5.7008f
C686 avss.n288 dvss 4.35256f
C687 avss.n289 dvss 2.30248f
C688 avss.n301 dvss 2.3148f
C689 avss.n302 dvss 4.37718f
C690 avss.n309 dvss 4.35256f
C691 avss.n310 dvss 2.17936f
C692 avss.n317 dvss 17.3824f
C693 avss.n356 dvss 1.80693f
C694 avss.n377 dvss 1.80693f
C695 avss.n418 dvss 1.80693f
C696 avss.n429 dvss 1.94342f
C697 avss.n431 dvss 1.94342f
C698 avss.n484 dvss 5.94779f
C699 avss.n485 dvss 6.68171f
C700 avss.n486 dvss 9.88291f
C701 avss.n487 dvss 4.16193f
C702 avss.n488 dvss 40.396103f
C703 avss.n489 dvss 26.021599f
C704 avss.n501 dvss 1.06406f
C705 avss.n557 dvss 1.94342f
C706 avss.n571 dvss 1.80693f
C707 avss.t152 dvss 7.01827f
C708 avss.n585 dvss 6.64036f
C709 avss.n591 dvss 4.83181f
C710 avss.n592 dvss 9.85383f
C711 avss.n593 dvss 3.43526f
C712 avss.t61 dvss 5.7008f
C713 avss.n602 dvss 2.05623f
C714 avss.n612 dvss 1.80693f
C715 avss.n623 dvss 1.94342f
C716 avss.n634 dvss 2.95744f
C717 avss.n635 dvss 5.89287f
C718 avss.n636 dvss 3.56744f
C719 avss.n637 dvss 2.61079f
C720 avss.t25 dvss 2.8988f
C721 avss.n647 dvss 4.16246f
C722 avss.n648 dvss 3.48605f
C723 avss.n654 dvss 2.48054f
C724 avss.n655 dvss 38.3629f
C725 avss.n656 dvss 33.1972f
C726 avss.n657 dvss 6.21863f
C727 avss.n658 dvss 6.23994f
C728 avss.n694 dvss 8.86258f
C729 avss.n705 dvss 1.18123f
C730 avss.n713 dvss 6.30083f
C731 avss.n719 dvss 3.95622f
C732 avss.n720 dvss 21.1607f
C733 avss.n721 dvss 6.11833f
C734 avss.n722 dvss 6.03898f
C735 avss.n723 dvss 5.55681f
C736 avss.n724 dvss 5.75446f
C737 avss.n725 dvss 1.45429f
C738 avss.n726 dvss 1.4843f
C739 avss.n727 dvss 1.79671f
C740 avss.t80 dvss 24.9958f
C741 avss.n731 dvss 1.84429f
C742 avss.n732 dvss 4.9089f
C743 avss.n733 dvss 6.53045f
C744 avss.n734 dvss 2.40661f
C745 avss.t10 dvss 86.8916f
C746 avss.n735 dvss 2.40661f
C747 avss.n736 dvss 24.0401f
C748 avss.n737 dvss 10.747499f
C749 avss.n738 dvss 13.144401f
C750 avss.n739 dvss 16.679f
C751 avss.n740 dvss 18.5431f
C752 multiplexer_0.vtrip_1.n0 dvss 1.46136f
C753 multiplexer_0.vtrip_1.n1 dvss 1.3392f
C754 multiplexer_0.vtrip_1.t12 dvss 1.05095f
C755 multiplexer_0.vtrip_1.n2 dvss 2.1732f
C756 multiplexer_0.vtrip_1.n3 dvss 1.85466f
C757 multiplexer_0.vtrip_1.t7 dvss 1.00152f
C758 multiplexer_0.vtrip_1.n4 dvss 1.93214f
C759 multiplexer_0.vtrip_1.n5 dvss 1.85466f
C760 multiplexer_0.vtrip_1.t3 dvss 1.00152f
C761 multiplexer_0.vtrip_1.n6 dvss 1.39736f
C762 multiplexer_0.vtrip_1.n7 dvss 1.85466f
C763 multiplexer_0.vtrip_1.t9 dvss 1.00152f
C764 multiplexer_0.vtrip_1.t8 dvss 1.0902f
C765 multiplexer_0.vtrip_1.n8 dvss 1.33919f
C766 multiplexer_0.vtrip_1.t6 dvss 1.05073f
C767 multiplexer_0.vtrip_1.n10 dvss 1.21589f
C768 multiplexer_0.vtrip_1.n11 dvss 3.1186f
.ends


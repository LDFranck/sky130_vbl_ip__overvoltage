magic
tech sky130A
timestamp 1712777902
<< pwell >>
rect -1098 -155 1098 155
<< nmos >>
rect -1000 -50 1000 50
<< ndiff >>
rect -1029 44 -1000 50
rect -1029 -44 -1023 44
rect -1006 -44 -1000 44
rect -1029 -50 -1000 -44
rect 1000 44 1029 50
rect 1000 -44 1006 44
rect 1023 -44 1029 44
rect 1000 -50 1029 -44
<< ndiffc >>
rect -1023 -44 -1006 44
rect 1006 -44 1023 44
<< psubdiff >>
rect -1080 120 -1032 137
rect 1032 120 1080 137
rect -1080 89 -1063 120
rect 1063 89 1080 120
rect -1080 -120 -1063 -89
rect 1063 -120 1080 -89
rect -1080 -137 -1032 -120
rect 1032 -137 1080 -120
<< psubdiffcont >>
rect -1032 120 1032 137
rect -1080 -89 -1063 89
rect 1063 -89 1080 89
rect -1032 -137 1032 -120
<< poly >>
rect -1000 86 1000 94
rect -1000 69 -992 86
rect 992 69 1000 86
rect -1000 50 1000 69
rect -1000 -69 1000 -50
rect -1000 -86 -992 -69
rect 992 -86 1000 -69
rect -1000 -94 1000 -86
<< polycont >>
rect -992 69 992 86
rect -992 -86 992 -69
<< locali >>
rect -1080 120 -1032 137
rect 1032 120 1080 137
rect -1080 89 -1063 120
rect 1063 89 1080 120
rect -1000 69 -992 86
rect 992 69 1000 86
rect -1023 44 -1006 52
rect -1023 -52 -1006 -44
rect 1006 44 1023 52
rect 1006 -52 1023 -44
rect -1000 -86 -992 -69
rect 992 -86 1000 -69
rect -1080 -120 -1063 -89
rect 1063 -120 1080 -89
rect -1080 -137 -1032 -120
rect 1032 -137 1080 -120
<< viali >>
rect -992 69 992 86
rect -1023 -44 -1006 44
rect 1006 -44 1023 44
rect -992 -86 992 -69
<< metal1 >>
rect -998 86 998 89
rect -998 69 -992 86
rect 992 69 998 86
rect -998 66 998 69
rect -1026 44 -1003 50
rect -1026 -44 -1023 44
rect -1006 -44 -1003 44
rect -1026 -50 -1003 -44
rect 1003 44 1026 50
rect 1003 -44 1006 44
rect 1023 -44 1026 44
rect 1003 -50 1026 -44
rect -998 -69 998 -66
rect -998 -86 -992 -69
rect 992 -86 998 -69
rect -998 -89 998 -86
<< properties >>
string FIXED_BBOX -1071 -128 1071 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 20.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

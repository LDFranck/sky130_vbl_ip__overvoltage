magic
tech sky130A
magscale 1 2
timestamp 1712755851
<< nwell >>
rect -496 -319 496 319
<< pmos >>
rect -300 -100 300 100
<< pdiff >>
rect -358 88 -300 100
rect -358 -88 -346 88
rect -312 -88 -300 88
rect -358 -100 -300 -88
rect 300 88 358 100
rect 300 -88 312 88
rect 346 -88 358 88
rect 300 -100 358 -88
<< pdiffc >>
rect -346 -88 -312 88
rect 312 -88 346 88
<< nsubdiff >>
rect -460 249 -364 283
rect 364 249 460 283
rect -460 187 -426 249
rect 426 187 460 249
rect -460 -249 -426 -187
rect 426 -249 460 -187
rect -460 -283 -364 -249
rect 364 -283 460 -249
<< nsubdiffcont >>
rect -364 249 364 283
rect -460 -187 -426 187
rect 426 -187 460 187
rect -364 -283 364 -249
<< poly >>
rect -300 181 300 197
rect -300 147 -284 181
rect 284 147 300 181
rect -300 100 300 147
rect -300 -147 300 -100
rect -300 -181 -284 -147
rect 284 -181 300 -147
rect -300 -197 300 -181
<< polycont >>
rect -284 147 284 181
rect -284 -181 284 -147
<< locali >>
rect -460 249 -364 283
rect 364 249 460 283
rect -460 187 -426 249
rect 426 187 460 249
rect -300 147 -284 181
rect 284 147 300 181
rect -346 88 -312 104
rect -346 -104 -312 -88
rect 312 88 346 104
rect 312 -104 346 -88
rect -300 -181 -284 -147
rect 284 -181 300 -147
rect -460 -249 -426 -187
rect 426 -249 460 -187
rect -460 -283 -364 -249
rect 364 -283 460 -249
<< viali >>
rect -284 147 284 181
rect -346 -88 -312 88
rect 312 -88 346 88
rect -284 -181 284 -147
<< metal1 >>
rect -296 181 296 187
rect -296 147 -284 181
rect 284 147 296 181
rect -296 141 296 147
rect -352 88 -306 100
rect -352 -88 -346 88
rect -312 -88 -306 88
rect -352 -100 -306 -88
rect 306 88 352 100
rect 306 -88 312 88
rect 346 -88 352 88
rect 306 -100 352 -88
rect -296 -147 296 -141
rect -296 -181 -284 -147
rect 284 -181 296 -147
rect -296 -187 296 -181
<< properties >>
string FIXED_BBOX -443 -266 443 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 3.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

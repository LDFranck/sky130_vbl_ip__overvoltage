* NGSPICE file created from toplevel.ext - technology: sky130A

.subckt sky130_fd_pr__res_xhigh_po_1p41_LV9PDH a_8742_125# a_n3732_n557# a_1560_125#
+ a_3828_n557# a_n7512_n557# a_804_n557# a_7608_n557# a_n4110_n557# a_3072_125# a_4206_n557#
+ a_4584_125# a_n4110_125# a_6096_125# a_n5622_125# a_6852_n557# a_n4866_n557# a_n1464_n557#
+ a_3450_n557# a_48_125# a_n8646_n557# a_7230_n557# a_n5244_n557# a_n7134_125# a_n8646_125#
+ a_n1464_125# a_n9024_n557# a_n2976_125# a_804_125# a_2316_125# a_3828_125# a_n7890_n557#
+ a_5340_125# a_7986_n557# a_n4488_125# a_4584_n557# a_n2598_n557# a_1182_n557# a_6852_125#
+ a_8364_n557# a_n6378_n557# a_8364_125# a_1182_125# a_2694_125# a_n2220_125# a_n1842_n557#
+ a_48_n557# a_1938_n557# a_n3732_125# a_n708_125# a_n5622_n557# a_n2220_n557# a_5718_n557#
+ a_2316_n557# a_6096_n557# a_n5244_125# a_n6000_n557# a_n6756_125# a_7608_125# a_n8268_125#
+ a_n2976_n557# a_4962_n557# a_n1086_125# a_1560_n557# a_1938_125# a_n2598_125# a_3450_125#
+ a_4962_125# a_8742_n557# a_5340_n557# a_n6756_n557# a_426_125# a_n3354_n557# a_6474_125#
+ a_n7134_n557# a_426_n557# a_7986_125# a_n708_n557# a_n6000_125# a_n7512_125# a_2694_n557#
+ a_n1842_125# a_6474_n557# a_3072_n557# a_n4488_n557# a_n1086_n557# a_n330_125# a_n9024_125#
+ a_n3354_125# a_n8268_n557# a_n4866_125# a_n330_n557# a_n7890_125# a_4206_125# a_5718_125#
+ a_7230_125# VSUBS a_n6378_125#
X0 a_n8646_125# a_n8646_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X1 a_n6000_125# a_n6000_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X2 a_n1464_125# a_n1464_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X3 a_6474_125# a_6474_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X4 a_804_125# a_804_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X5 a_n7134_125# a_n7134_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X6 a_n4488_125# a_n4488_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X7 a_5718_125# a_5718_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X8 a_n1842_125# a_n1842_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X9 a_6852_125# a_6852_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X10 a_n7512_125# a_n7512_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X11 a_n4866_125# a_n4866_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X12 a_4206_125# a_4206_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X13 a_5340_125# a_5340_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X14 a_n330_125# a_n330_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X15 a_2694_125# a_2694_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X16 a_n7890_125# a_n7890_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X17 a_n3354_125# a_n3354_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X18 a_n2220_125# a_n2220_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X19 a_8364_125# a_8364_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X20 a_1182_125# a_1182_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X21 a_1938_125# a_1938_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X22 a_n9024_125# a_n9024_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X23 a_n708_125# a_n708_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X24 a_48_125# a_48_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X25 a_n6378_125# a_n6378_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X26 a_n3732_125# a_n3732_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X27 a_7608_125# a_7608_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X28 a_8742_125# a_8742_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X29 a_1560_125# a_1560_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X30 a_n6756_125# a_n6756_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X31 a_7230_125# a_7230_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X32 a_4584_125# a_4584_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X33 a_n5244_125# a_n5244_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X34 a_n4110_125# a_n4110_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X35 a_n2598_125# a_n2598_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X36 a_3072_125# a_3072_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X37 a_3828_125# a_3828_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X38 a_4962_125# a_4962_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X39 a_n8268_125# a_n8268_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X40 a_n5622_125# a_n5622_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X41 a_n2976_125# a_n2976_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X42 a_n1086_125# a_n1086_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X43 a_6096_125# a_6096_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X44 a_7986_125# a_7986_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X45 a_426_125# a_426_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X46 a_2316_125# a_2316_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
X47 a_3450_125# a_3450_n557# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=1.41
.ends

.subckt sky130_fd_pr__res_xhigh_po_1p41_H3F4MM a_1182_1930# a_n4488_n1826# a_7986_n1826#
+ a_n6378_n2362# a_n7890_5150# a_n7890_n5582# a_7986_5150# a_4584_5150# a_n2598_5150#
+ a_1182_5150# a_8364_1930# a_n6378_1930# a_n4866_n1826# a_n6756_n2362# a_8364_5150#
+ a_n6378_5150# a_n2598_n1826# a_n6000_n5582# a_n4488_n2362# a_n3732_1394# a_7986_n2362#
+ a_3828_1394# a_426_n5582# a_7230_n5582# a_7608_n5582# a_n2976_n1826# a_n4866_n2362#
+ a_n7512_1394# a_n4110_1394# a_804_1394# a_7608_1394# a_4206_1394# a_4206_n1826#
+ a_n1842_1930# a_n4110_n5582# a_804_n5582# a_n2598_n2362# a_48_1930# a_1938_1930#
+ a_5340_n5582# a_n1842_5150# a_5718_n5582# a_48_5150# a_1938_5150# a_n5622_1930#
+ a_n2976_n2362# a_n2220_1930# a_5718_1930# a_3072_n5582# a_2316_1930# a_n9024_n1826#
+ a_6096_1930# a_2316_n1826# a_4206_n2362# a_n2220_n5582# a_n5622_5150# a_n2220_5150#
+ a_5718_5150# a_2316_5150# a_6852_1394# a_n6000_1930# a_6096_5150# a_n4866_1394#
+ a_3450_1394# a_3450_n5582# a_3828_n5582# a_n1464_1394# a_n8268_n5582# a_n6000_5150#
+ a_1182_n5582# a_n7134_n1826# a_n9024_n2362# a_2316_n2362# a_n8646_1394# a_7230_1394#
+ a_n5244_1394# a_8364_n1826# a_4962_1930# a_n2976_1930# a_1560_1930# a_n8646_n5582#
+ a_1560_n5582# a_n7512_n1826# a_1938_n5582# a_6096_n1826# a_n9024_1394# a_4962_5150#
+ a_n2976_5150# a_n6378_n5582# a_n5244_n1826# a_n7134_n2362# a_1560_5150# a_8742_n1826#
+ a_8742_1930# a_n6756_1930# a_5340_1930# a_n3354_1930# a_n330_n1826# a_6474_n1826#
+ a_n708_n1826# a_8364_n2362# a_8742_5150# a_n6756_n5582# a_n6756_5150# a_n5622_n1826#
+ a_5340_5150# a_n7512_n2362# a_48_n1826# a_n7890_1394# a_n3354_5150# a_6096_n2362#
+ a_n7134_1930# a_7986_1394# a_n4488_n5582# a_426_1930# a_4584_1394# a_7986_n5582#
+ a_n3354_n1826# a_n2598_1394# a_6852_n1826# a_n5244_n2362# a_8742_n2362# a_1182_1394#
+ a_n708_1930# a_n7134_5150# a_n1086_n1826# a_426_5150# a_4584_n1826# a_n330_n2362#
+ a_6474_n2362# a_n708_n2362# a_8364_1394# a_n4866_n5582# a_n3732_n1826# a_n6378_1394#
+ a_n5622_n2362# a_48_n2362# a_n708_5150# a_2694_1930# a_n2598_n5582# a_n1464_n1826#
+ a_4962_n1826# a_n3354_n2362# a_6852_n2362# a_2694_5150# a_2694_n1826# a_n1086_n2362#
+ a_4584_n2362# a_6474_1930# a_n2976_n5582# a_n4488_1930# a_n1842_n1826# a_n3732_n2362#
+ a_3072_1930# a_n1086_1930# a_4206_n5582# a_6474_5150# a_n1464_n2362# a_4962_n2362#
+ a_n4488_5150# a_3072_5150# a_n1842_1394# a_n1086_5150# a_n8268_1930# a_48_1394#
+ a_1938_1394# a_2694_n2362# a_n330_1930# a_n1842_n2362# a_n8268_5150# a_n5622_1394#
+ a_n9024_n5582# a_n2220_1394# a_2316_n5582# a_5718_1394# a_n7890_n1826# a_n330_5150#
+ a_2316_1394# a_6096_1394# a_n6000_1394# a_n3732_1930# a_n7134_n5582# a_3828_1930#
+ a_n6000_n1826# a_n7890_n2362# a_n3732_5150# a_8364_n5582# a_426_n1826# a_7230_n1826#
+ a_3828_5150# a_7608_n1826# a_n7512_1930# a_n7512_n5582# a_n4110_1930# a_804_1930#
+ a_7608_1930# a_4962_1394# a_n2976_1394# a_4206_1930# a_1560_1394# a_6096_n5582#
+ a_n7512_5150# a_n5244_n5582# a_n4110_n1826# a_8742_n5582# a_804_n1826# a_n6000_n2362#
+ a_n4110_5150# a_804_5150# a_7608_5150# a_4206_5150# a_8742_1394# a_n6756_1394# a_5340_1394#
+ a_n3354_1394# a_6474_n5582# a_n330_n5582# a_n708_n5582# a_5340_n1826# a_426_n2362#
+ a_5718_n1826# a_7230_n2362# a_7608_n2362# a_n5622_n5582# a_48_n5582# a_3072_n1826#
+ a_n7134_1394# a_n3354_n5582# a_6852_n5582# a_n2220_n1826# a_n4110_n2362# a_804_n2362#
+ a_426_1394# a_6852_1930# a_n4866_1930# a_3450_1930# a_n1464_1930# a_n1086_n5582#
+ a_4584_n5582# a_n708_1394# a_3450_n1826# a_5340_n2362# a_3828_n1826# a_5718_n2362#
+ a_n3732_n5582# a_6852_5150# a_n4866_5150# a_3450_5150# a_n1464_5150# a_n8268_n1826#
+ a_1182_n1826# a_n8646_1930# a_3072_n2362# a_7230_1930# a_n5244_1930# a_n1464_n5582#
+ a_4962_n5582# a_n2220_n2362# a_2694_1394# a_n8646_5150# a_7230_5150# a_2694_n5582#
+ a_n8646_n1826# a_n5244_5150# a_1560_n1826# a_1938_n1826# a_3450_n2362# a_3828_n2362#
+ a_n9024_1930# a_n1842_n5582# a_6474_1394# a_n4488_1394# a_3072_1394# a_n6378_n1826#
+ a_n8268_n2362# a_n1086_1394# a_1182_n2362# a_n9024_5150# a_n8268_1394# a_n7890_1930#
+ a_n6756_n1826# a_n8646_n2362# a_1560_n2362# a_1938_n2362# a_7986_1930# VSUBS a_4584_1930#
+ a_n2598_1930# a_n330_1394#
X0 a_n1464_n2362# a_n1464_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X1 a_n3732_n2362# a_n3732_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X2 a_426_n2362# a_426_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X3 a_n4110_5150# a_n4110_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X4 a_n5244_5150# a_n5244_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X5 a_n2598_5150# a_n2598_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X6 a_3072_5150# a_3072_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X7 a_3828_5150# a_3828_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X8 a_4962_5150# a_4962_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X9 a_n9024_1394# a_n9024_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X10 a_6474_1394# a_6474_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X11 a_n8268_5150# a_n8268_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X12 a_8742_1394# a_8742_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X13 a_5718_1394# a_5718_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X14 a_n330_1394# a_n330_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X15 a_n9024_n2362# a_n9024_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X16 a_3072_1394# a_3072_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X17 a_n7890_1394# a_n7890_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X18 a_n5622_5150# a_n5622_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X19 a_5340_1394# a_5340_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X20 a_2316_1394# a_2316_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X21 a_n1086_5150# a_n1086_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X22 a_6096_5150# a_6096_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X23 a_6474_n2362# a_6474_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X24 a_8742_n2362# a_8742_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X25 a_5718_n2362# a_5718_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X26 a_n330_n2362# a_n330_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X27 a_7986_5150# a_7986_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X28 a_n4488_1394# a_n4488_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X29 a_n2976_5150# a_n2976_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X30 a_2316_5150# a_2316_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X31 a_n6756_1394# a_n6756_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X32 a_426_5150# a_426_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X33 a_3450_5150# a_3450_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X34 a_3072_n2362# a_3072_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X35 a_n7890_n2362# a_n7890_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X36 a_5340_n2362# a_5340_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X37 a_2316_n2362# a_2316_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X38 a_n1086_1394# a_n1086_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X39 a_n3354_1394# a_n3354_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X40 a_n4488_n2362# a_n4488_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X41 a_n5622_1394# a_n5622_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X42 a_n6756_n2362# a_n6756_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X43 a_n1086_n2362# a_n1086_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X44 a_n8646_5150# a_n8646_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X45 a_n3354_n2362# a_n3354_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X46 a_n5622_n2362# a_n5622_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X47 a_n6000_5150# a_n6000_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X48 a_6474_5150# a_6474_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X49 a_n1464_5150# a_n1464_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X50 a_804_5150# a_804_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X51 a_n7134_5150# a_n7134_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X52 a_6096_1394# a_6096_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X53 a_n4488_5150# a_n4488_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X54 a_8364_1394# a_8364_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X55 a_7608_1394# a_7608_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X56 a_n1842_5150# a_n1842_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X57 a_5718_5150# a_5718_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X58 a_6852_5150# a_6852_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X59 a_6096_n2362# a_6096_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X60 a_7230_1394# a_7230_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X61 a_4206_1394# a_4206_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X62 a_8364_n2362# a_8364_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X63 a_7608_n2362# a_7608_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X64 a_n6378_1394# a_n6378_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X65 a_n8646_1394# a_n8646_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X66 a_7230_n2362# a_7230_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X67 a_4206_n2362# a_4206_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X68 a_n2220_1394# a_n2220_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X69 a_n5244_1394# a_n5244_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X70 a_n6378_n2362# a_n6378_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X71 a_n7512_1394# a_n7512_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X72 a_n7512_5150# a_n7512_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X73 a_n8646_n2362# a_n8646_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X74 a_2694_1394# a_2694_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X75 a_n4866_5150# a_n4866_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X76 a_4206_5150# a_4206_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X77 a_4962_1394# a_4962_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X78 a_1938_1394# a_1938_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X79 a_5340_5150# a_5340_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X80 a_n2220_n2362# a_n2220_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X81 a_n5244_n2362# a_n5244_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X82 a_n7512_n2362# a_n7512_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X83 a_n330_5150# a_n330_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X84 a_2694_5150# a_2694_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X85 a_1560_1394# a_1560_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X86 a_2694_n2362# a_2694_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X87 a_4962_n2362# a_4962_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X88 a_1938_n2362# a_1938_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X89 a_48_1394# a_48_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X90 a_n2976_1394# a_n2976_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X91 a_1560_n2362# a_1560_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X92 a_48_n2362# a_48_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X93 a_n7890_5150# a_n7890_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X94 a_n1842_1394# a_n1842_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X95 a_n2220_5150# a_n2220_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X96 a_n2976_n2362# a_n2976_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X97 a_n3354_5150# a_n3354_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X98 a_8364_5150# a_8364_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X99 a_804_1394# a_804_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X100 a_1182_5150# a_1182_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X101 a_n1842_n2362# a_n1842_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X102 a_1938_5150# a_1938_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X103 a_804_n2362# a_804_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X104 a_n708_5150# a_n708_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X105 a_48_5150# a_48_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X106 a_n9024_5150# a_n9024_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X107 a_n8268_1394# a_n8268_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X108 a_n6378_5150# a_n6378_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X109 a_n3732_5150# a_n3732_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X110 a_7608_5150# a_7608_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X111 a_8742_5150# a_8742_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X112 a_7986_1394# a_7986_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X113 a_n4110_1394# a_n4110_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X114 a_n7134_1394# a_n7134_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X115 a_n8268_n2362# a_n8268_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X116 a_4584_1394# a_4584_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X117 a_1560_5150# a_1560_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X118 a_6852_1394# a_6852_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X119 a_3828_1394# a_3828_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X120 a_7986_n2362# a_7986_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X121 a_n4110_n2362# a_n4110_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X122 a_n7134_n2362# a_n7134_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X123 a_n708_1394# a_n708_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X124 a_1182_1394# a_1182_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X125 a_n6000_1394# a_n6000_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X126 a_3450_1394# a_3450_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X127 a_4584_n2362# a_4584_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X128 a_6852_n2362# a_6852_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X129 a_3828_n2362# a_3828_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X130 a_n2598_1394# a_n2598_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X131 a_n708_n2362# a_n708_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X132 a_n4866_1394# a_n4866_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X133 a_n6756_5150# a_n6756_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X134 a_1182_n2362# a_1182_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X135 a_n6000_n2362# a_n6000_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X136 a_7230_5150# a_7230_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X137 a_3450_n2362# a_3450_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X138 a_n1464_1394# a_n1464_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X139 a_4584_5150# a_4584_1930# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X140 a_n2598_n2362# a_n2598_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X141 a_n3732_1394# a_n3732_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X142 a_n4866_n2362# a_n4866_n5582# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
X143 a_426_1394# a_426_n1826# VSUBS sky130_fd_pr__res_xhigh_po_1p41 l=14.1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8 a_300_n300# a_n492_n522# a_n358_n300#
+ a_n300_n388#
X0 a_300_n300# a_n300_n388# a_n358_n300# a_n492_n522# sky130_fd_pr__nfet_g5v0d10v5 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=3
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_F6RBXN a_n147_n172# a_n45_n70#
D0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 pj=2.3e+06 area=3.15e+11
.ends

.subckt voltage_divider out_0000 out_0001 out_0010 out_0011 out_0100 out_0101 out_0110
+ out_0111 out_1000 out_1001 out_1010 out_1011 out_1100 out_1101 out_1110 out_1111
+ ena avdd avss
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_0 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_LV9PDH_2 avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss avss
+ avss avss avss avss avss avss avss avss avss sky130_fd_pr__res_xhigh_po_1p41_LV9PDH
Xsky130_fd_pr__res_xhigh_po_1p41_H3F4MM_0 m1_3399_9649# m1_7155_3979# m1_7155_16831#
+ m1_7155_2467# m1_179_955# m1_10911_577# m1_179_16831# m1_179_13051# m1_179_6247#
+ m1_179_10027# m1_3399_17209# m1_3399_2467# m1_7155_3979# m1_7155_2089# m1_179_16831#
+ m1_179_2467# m1_7155_6247# m1_10911_2845# out_1110 m1_3935_5113# m1_7155_16831#
+ m1_3935_12673# out_0011 m1_10911_15697# m1_10911_16453# m1_7155_5491# out_1110 m1_3399_1333#
+ m1_3935_4357# m1_3935_9649# m1_3935_16453# m1_3935_12673# m1_7155_13051# m1_3399_6625#
+ out_1101 out_0010 out_1000 m1_3399_8893# m1_3399_10405# m1_10911_14185# m1_179_7003#
+ m1_10911_14185# m1_179_8515# m1_179_10783# m1_3399_3223# out_1010 m1_3399_6625#
+ m1_3399_14185# m1_10911_11917# m1_3399_11161# avss m1_3399_14941# m1_7155_10783#
+ m1_7691_13051# out_0111 m1_179_3223# m1_179_6247# m1_179_14563# m1_179_10783# m1_3935_15697#
+ m1_3399_2845# m1_179_14563# m1_3399_3979# m1_3935_11917# m1_10911_11917# m1_10911_12673#
+ m1_3935_7381# m1_10911_577# m1_179_2467# out_0010 m1_7155_1711# avss m1_7691_10783#
+ m1_3399_199# m1_3935_15697# m1_3399_3601# m1_7155_17209# m1_3399_13429# m1_3399_5869#
+ m1_3399_10405# m1_10901_199# out_0001 m1_7155_1333# out_0001 m1_7155_14563# avss
+ m1_179_13807# m1_179_5491# m1_10911_2089# m1_7155_3601# m1_7155_1711# m1_179_10027#
+ avss avss m1_3399_2089# m1_3399_14185# m1_3399_5113# m1_7155_8515# m1_7155_15319#
+ m1_7155_7759# m1_7155_17209# avss m1_10911_2089# m1_179_1711# m1_7155_3223# m1_179_13807#
+ m1_7155_1333# m1_7155_8515# m1_3399_955# m1_179_5491# m1_7691_14563# m1_3399_1711#
+ m1_3935_16453# out_1101 m1_3399_8893# m1_3935_13429# m1_10911_16453# m1_7155_5491#
+ m1_3935_5869# m1_7155_15319# m1_7155_3601# avss m1_3935_9649# m1_3399_8137# m1_179_1711#
+ m1_7155_7759# m1_179_9271# m1_7155_13051# out_0100 m1_7691_15319# out_0101 m1_3399_17209#
+ out_1111 m1_7155_4735# m1_3399_2467# m1_7155_3223# out_0100 m1_179_7759# m1_3399_11161#
+ out_1001 m1_7155_7003# m1_7155_13807# out_1010 m1_7691_15319# m1_179_11539# m1_7155_11539#
+ out_0101 m1_7691_13051# m1_3399_14941# out_1001 m1_3399_4357# m1_7155_7003# out_1100
+ m1_3399_11917# m1_3399_7381# m1_10911_12673# m1_179_15319# m1_7691_7003# m1_7691_13807#
+ m1_179_3979# m1_179_11539# m1_3935_6625# m1_179_7759# m1_3399_577# m1_3935_8893#
+ m1_3935_10405# 51 m1_3399_8137# m1_7691_7003# m1_179_199# m1_3399_3223# avss m1_3935_6625#
+ out_0000 m1_3935_14185# m1_7155_955# m1_179_8515# m1_3935_11161# m1_3935_14941#
+ m1_3399_2845# m1_3399_5113# m1_10911_1333# m1_3399_12673# m1_7155_2845# m1_7155_955#
+ m1_179_4735# avdd m1_7155_9271# m1_7155_16075# m1_179_12295# m1_7155_16075# m1_3399_1333#
+ m1_10911_1333# m1_3399_4357# m1_3399_9649# m1_3399_16453# m1_3935_13429# m1_3935_5869#
+ m1_3399_12673# m1_3935_10405# m1_10911_14941# m1_179_955# out_1111 m1_7155_4735#
+ avss m1_7155_9271# m1_7155_2845# m1_179_4735# m1_179_9271# m1_179_16075# m1_179_13051#
+ avss m1_3399_2089# m1_3935_14185# m1_3935_5113# m1_10911_14941# m1_10901_8137# m1_10901_8137#
+ m1_7155_13807# m1_7691_9271# m1_7155_14563# m1_7691_16075# m1_7691_16075# m1_10911_2845#
+ out_0011 m1_7155_11539# m1_3399_1711# out_1011 m1_10911_15697# m1_7155_6247# out_1100
+ m1_7691_9271# m1_3935_8893# m1_3399_15697# m1_3399_3979# m1_3399_11917# m1_3399_7381#
+ out_0110 m1_10911_13429# m1_3935_8137# m1_7155_12295# m1_7691_13807# m1_7155_12295#
+ m1_7691_14563# out_1011 m1_179_15319# m1_179_3979# m1_179_12295# m1_179_7003# m1_7155_577#
+ m1_7155_10027# m1_3399_199# 51 m1_3399_15697# m1_3399_3601# out_0110 m1_10911_13429#
+ out_1000 m1_3935_11161# m1_179_199# m1_179_16075# out_0000 m1_7155_199# m1_179_3223#
+ m1_7155_10027# m1_7155_10783# m1_7691_12295# m1_7691_12295# avss out_0111 m1_3935_14941#
+ m1_3935_4357# m1_3935_11917# m1_7155_2467# m1_7155_577# m1_3935_7381# m1_7691_10027#
+ avss m1_3399_577# m1_3399_955# m1_7155_2089# m1_7155_199# m1_7691_10027# m1_7691_10783#
+ m1_3399_16453# avss m1_3399_13429# m1_3399_5869# m1_3935_8137# sky130_fd_pr__res_xhigh_po_1p41_H3F4MM
Xsky130_fd_pr__nfet_g5v0d10v5_SB5CJ8_0 avss avss m1_10901_199# ena sky130_fd_pr__nfet_g5v0d10v5_SB5CJ8
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 avss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CY564Z a_300_n100# a_n492_n322# a_n358_n100#
+ a_n300_n188#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n492_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt trans_gate_m in ena_b ena out avdd vss
Xsky130_fd_pr__pfet_g5v0d10v5_6H9SQ3_1 ena_b out avdd in sky130_fd_pr__pfet_g5v0d10v5_6H9SQ3
Xsky130_fd_pr__nfet_g5v0d10v5_CY564Z_0 out vss in ena sky130_fd_pr__nfet_g5v0d10v5_CY564Z
.ends

.subckt multiplexer in_0000 in_0001 in_0010 in_0011 in_0100 in_0101 in_0110 in_0111
+ vtrip_3 vtrip_3_b vtrip_2 vtrip_1 out vtrip_1_b vtrip_0 in_1000 in_1001 in_1010
+ in_1011 in_1100 in_1101 in_1110 in_1111 vtrip_2_b vtrip_0_b vss avdd
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_3 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_2 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_4 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_5 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_6 vss vtrip_1_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_7 vss vtrip_1 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_8 vss vtrip_2_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_9 vss vtrip_2 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_31 trans_gate_m_31/in vtrip_1 vtrip_1_b trans_gate_m_20/in avdd vss
+ trans_gate_m
Xtrans_gate_m_20 trans_gate_m_20/in vtrip_2 vtrip_2_b trans_gate_m_33/in avdd vss
+ trans_gate_m
Xtrans_gate_m_0 in_0010 vtrip_0 vtrip_0_b trans_gate_m_29/in avdd vss trans_gate_m
Xtrans_gate_m_1 in_0011 vtrip_0_b vtrip_0 trans_gate_m_29/in avdd vss trans_gate_m
Xtrans_gate_m_32 trans_gate_m_32/in vtrip_2 vtrip_2_b trans_gate_m_34/in avdd vss
+ trans_gate_m
Xtrans_gate_m_10 in_1000 vtrip_0 vtrip_0_b trans_gate_m_23/in avdd vss trans_gate_m
Xtrans_gate_m_21 trans_gate_m_5/out vtrip_1_b vtrip_1 trans_gate_m_32/in avdd vss
+ trans_gate_m
Xtrans_gate_m_2 in_0110 vtrip_0 vtrip_0_b trans_gate_m_3/out avdd vss trans_gate_m
Xtrans_gate_m_33 trans_gate_m_33/in vtrip_3 vtrip_3_b out avdd vss trans_gate_m
Xtrans_gate_m_11 in_1001 vtrip_0_b vtrip_0 trans_gate_m_23/in avdd vss trans_gate_m
Xtrans_gate_m_3 in_0111 vtrip_0_b vtrip_0 trans_gate_m_3/out avdd vss trans_gate_m
Xtrans_gate_m_12 in_0101 vtrip_0_b vtrip_0 trans_gate_m_27/in avdd vss trans_gate_m
Xtrans_gate_m_34 trans_gate_m_34/in vtrip_3_b vtrip_3 out avdd vss trans_gate_m
Xtrans_gate_m_23 trans_gate_m_23/in vtrip_1 vtrip_1_b trans_gate_m_32/in avdd vss
+ trans_gate_m
Xtrans_gate_m_13 in_0100 vtrip_0 vtrip_0_b trans_gate_m_27/in avdd vss trans_gate_m
Xtrans_gate_m_4 in_1011 vtrip_0_b vtrip_0 trans_gate_m_5/out avdd vss trans_gate_m
Xtrans_gate_m_14 in_0001 vtrip_0_b vtrip_0 trans_gate_m_31/in avdd vss trans_gate_m
Xtrans_gate_m_25 trans_gate_m_3/out vtrip_1_b vtrip_1 trans_gate_m_28/in avdd vss
+ trans_gate_m
Xtrans_gate_m_5 in_1010 vtrip_0 vtrip_0_b trans_gate_m_5/out avdd vss trans_gate_m
Xtrans_gate_m_15 in_0000 vtrip_0 vtrip_0_b trans_gate_m_31/in avdd vss trans_gate_m
Xtrans_gate_m_27 trans_gate_m_27/in vtrip_1 vtrip_1_b trans_gate_m_28/in avdd vss
+ trans_gate_m
Xtrans_gate_m_37 trans_gate_m_37/in vtrip_2_b vtrip_2 trans_gate_m_34/in avdd vss
+ trans_gate_m
Xtrans_gate_m_6 in_1110 vtrip_0 vtrip_0_b trans_gate_m_7/out avdd vss trans_gate_m
Xtrans_gate_m_28 trans_gate_m_28/in vtrip_2_b vtrip_2 trans_gate_m_33/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_10 vss vtrip_3_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_7 in_1111 vtrip_0_b vtrip_0 trans_gate_m_7/out avdd vss trans_gate_m
Xtrans_gate_m_29 trans_gate_m_29/in vtrip_1_b vtrip_1 trans_gate_m_20/in avdd vss
+ trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_11 vss vtrip_3 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xtrans_gate_m_18 trans_gate_m_9/out vtrip_1 vtrip_1_b trans_gate_m_37/in avdd vss
+ trans_gate_m
Xtrans_gate_m_8 in_1101 vtrip_0_b vtrip_0 trans_gate_m_9/out avdd vss trans_gate_m
Xtrans_gate_m_19 trans_gate_m_7/out vtrip_1_b vtrip_1 trans_gate_m_37/in avdd vss
+ trans_gate_m
Xtrans_gate_m_9 in_1100 vtrip_0 vtrip_0_b trans_gate_m_9/out avdd vss trans_gate_m
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 vss vtrip_0 sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_1 vss vtrip_0_b sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_YHAZV5 a_n300_n197# a_300_n100# w_n558_n397#
+ a_n358_n100#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n558_n397# sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__diode_pw2nd_05v5_37RBXE a_n147_n172# a_n45_n70#
D0 a_n147_n172# a_n45_n70# sky130_fd_pr__diode_pw2nd_05v5 pj=2.3e+06 area=3.15e+11
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_EEVBR7 a_n300_n288# a_300_n200# a_n492_n422#
+ a_n358_n200#
X0 a_300_n200# a_n300_n288# a_n358_n200# a_n492_n422# sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=3
.ends

.subckt sky130_fd_pr__nfet_01v8_MG6U6H a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9Q3 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt level_shifter in out out_b dvss avss li_5238_n1104# avdd
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0 out_b out avdd avdd sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1 out out_b avdd avdd sky130_fd_pr__pfet_g5v0d10v5_YHAZV5
Xsky130_fd_pr__diode_pw2nd_05v5_37RBXE_0 dvss in sky130_fd_pr__diode_pw2nd_05v5_37RBXE
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0 in_b out avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1 in out_b avss avss sky130_fd_pr__nfet_g5v0d10v5_EEVBR7
Xsky130_fd_pr__nfet_01v8_MG6U6H_0 dvss in_b in dvss sky130_fd_pr__nfet_01v8_MG6U6H
Xsky130_fd_pr__pfet_01v8_J2L9Q3_0 in in_b li_5238_n1104# li_5238_n1104# sky130_fd_pr__pfet_01v8_J2L9Q3
.ends

.subckt sky130_fd_pr__pfet_01v8_XTWSDC a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
.ends

.subckt sky130_fd_pr__nfet_01v8_7ZF23Z a_2000_n100# a_n2058_n100# a_n2000_n188# a_n2160_n274#
X0 a_2000_n100# a_n2000_n188# a_n2058_n100# a_n2160_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=20
.ends

.subckt sky130_fd_pr__nfet_01v8_V433WY a_300_n100# a_n358_n100# a_n300_n188# a_n460_n274#
X0 a_300_n100# a_n300_n188# a_n358_n100# a_n460_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_69BJMM a_n500_n188# a_500_n100# a_n692_n322#
+ a_n558_n100#
X0 a_500_n100# a_n500_n188# a_n558_n100# a_n692_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=5
.ends

.subckt sky130_fd_pr__pfet_g5v0d10v5_E7V9VM w_n758_n897# a_n558_n600# a_n500_n697#
+ a_500_n600#
X0 a_500_n600# a_n500_n697# a_n558_n600# w_n758_n897# sky130_fd_pr__pfet_g5v0d10v5 ad=1.74 pd=12.58 as=1.74 ps=12.58 w=6 l=5
.ends

.subckt trans_gate in ena_b ena out vss avdd
XXM1 ena out vss in sky130_fd_pr__nfet_g5v0d10v5_69BJMM
XXM2 avdd out ena_b in sky130_fd_pr__pfet_g5v0d10v5_E7V9VM
.ends

.subckt sky130_fd_pr__pfet_01v8_C2YSV5 a_n300_n197# a_300_n100# a_n358_n100# w_n496_n319#
X0 a_300_n100# a_n300_n197# a_n358_n100# w_n496_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=3
.ends

.subckt sky130_fd_pr__pfet_01v8_J2L9E5 w_n296_n319# a_n100_n197# a_100_n100# a_n158_n100#
X0 a_100_n100# a_n100_n197# a_n158_n100# w_n296_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_GGMWVD w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_CDT3CS a_n1600_n197# a_1600_n100# a_n1658_n100# w_n1796_n319#
X0 a_1600_n100# a_n1600_n197# a_n1658_n100# w_n1796_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=16
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z a_100_n100# a_n292_n322# a_n158_n100#
+ a_n100_n188#
X0 a_100_n100# a_n100_n188# a_n158_n100# a_n292_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=1
.ends

.subckt sky130_fd_pr__pfet_01v8_3HBZVM a_n158_n300# w_n296_n519# a_n100_n397# a_100_n300#
X0 a_100_n300# a_n100_n397# a_n158_n300# w_n296_n519# sky130_fd_pr__pfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt sky130_fd_pr__nfet_01v8_697RXD a_800_n100# a_n858_n100# a_n800_n188# a_n960_n274#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n960_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_4T6WVE a_100_n130# a_n292_n352# a_n158_n130#
+ a_n100_n218#
X0 a_100_n130# a_n100_n218# a_n158_n130# a_n292_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=1
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_6975WM a_800_n130# a_n992_n352# a_n858_n130#
+ a_n800_n218#
X0 a_800_n130# a_n800_n218# a_n858_n130# a_n992_n352# sky130_fd_pr__nfet_g5v0d10v5 ad=0.377 pd=3.18 as=0.377 ps=3.18 w=1.3 l=8
.ends

.subckt sky130_fd_pr__nfet_g5v0d10v5_DEN7YK a_800_n100# a_n992_n322# a_n858_n100#
+ a_n800_n188#
X0 a_800_n100# a_n800_n188# a_n858_n100# a_n992_n322# sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__pfet_01v8_G3L97A w_n996_n319# a_n800_n197# a_800_n100# a_n858_n100#
X0 a_800_n100# a_n800_n197# a_n858_n100# w_n996_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=8
.ends

.subckt sky130_fd_pr__nfet_01v8_C8TQ3N a_n158_n300# a_n100_n388# a_n260_n474# a_100_n300#
X0 a_100_n300# a_n100_n388# a_n158_n300# a_n260_n474# sky130_fd_pr__nfet_01v8 ad=0.87 pd=6.58 as=0.87 ps=6.58 w=3 l=1
.ends

.subckt comp_hyst out vref vin ena ibias dvss dvdd
XXMD16[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM12 dvss net1 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
XXM14 dvss net2 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXM13 dvss net5 ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
Xx1 ibias ena_b ena net5 dvss dvdd trans_gate
XXM15 ena net4 dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXM16 ena net3 dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXM17 dvss out ena_b dvss sky130_fd_pr__nfet_01v8_V433WY
XXMD1[19] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM18 ena ena_b dvdd dvdd sky130_fd_pr__pfet_01v8_C2YSV5
XXMD1[18] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM19 dvss ena_b ena dvss sky130_fd_pr__nfet_01v8_V433WY
XXM6[3] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM3[1] dvdd net4 net4 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[17] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[2] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXM3[0] dvdd net4 net4 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD1[16] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM6[1] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM6[0] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXMD1[15] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[13] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[14] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[9] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[12] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[8] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[11] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[7] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[10] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMDN1[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z
XXMD1[6] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXMD1[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XD1 dvss vref sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM7 dvdd net4 net2 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XD3 dvss ena sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXMD1[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM9 dvdd dvdd net3 out sky130_fd_pr__pfet_01v8_3HBZVM
XXM8 dvss net2 net2 dvss sky130_fd_pr__nfet_01v8_697RXD
XXMDN13[7] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXM1[1] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXMD1[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM1[0] net1 dvss net4 vref sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM4[1] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMDN13[6] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMD1[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_J2L9E5
XXM4[0] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8_CDT3CS
XXMDN13[5] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[4] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[3] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[2] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN13[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_4T6WVE
XXMDN8[1] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMDN8[0] dvss dvss dvss dvss sky130_fd_pr__nfet_g5v0d10v5_DEN7YK
XXMD16[5] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMD16[4] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[1] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[1] dvdd net4 net3 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[3] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM2[0] net1 dvss net3 vin sky130_fd_pr__nfet_g5v0d10v5_6975WM
XXM5[0] dvdd net4 net3 dvdd sky130_fd_pr__pfet_01v8_GGMWVD
XXMD16[2] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXMD8[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_G3L97A
Xsky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0 dvss vin sky130_fd_pr__diode_pw2nd_05v5_F6RBXN
XXM10 out net2 dvss dvss sky130_fd_pr__nfet_01v8_C8TQ3N
XXMD8[0] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_G3L97A
XXMD16[1] dvdd dvdd dvdd dvdd sky130_fd_pr__pfet_01v8_XTWSDC
XXM11 dvss net5 net5 dvss sky130_fd_pr__nfet_01v8_7ZF23Z
.ends

.subckt toplevel vtrip[3] vtrip[2] vtrip[1] vtrip[0] vbg ibias avdd dvss ena avss
+ dvdd ovout
Xvoltage_divider_0 multiplexer_0/in_0000 multiplexer_0/in_0001 multiplexer_0/in_0010
+ multiplexer_0/in_0011 multiplexer_0/in_0100 multiplexer_0/in_0101 multiplexer_0/in_0110
+ multiplexer_0/in_0111 multiplexer_0/in_1000 multiplexer_0/in_1001 multiplexer_0/in_1010
+ multiplexer_0/in_1011 multiplexer_0/in_1100 multiplexer_0/in_1101 multiplexer_0/in_1110
+ multiplexer_0/in_1111 ena avdd avss voltage_divider
Xmultiplexer_0 multiplexer_0/in_0000 multiplexer_0/in_0001 multiplexer_0/in_0010 multiplexer_0/in_0011
+ multiplexer_0/in_0100 multiplexer_0/in_0101 multiplexer_0/in_0110 multiplexer_0/in_0111
+ level_shifter_3/out level_shifter_3/out_b level_shifter_2/out level_shifter_1/out
+ vin level_shifter_1/out_b level_shifter_0/out multiplexer_0/in_1000 multiplexer_0/in_1001
+ multiplexer_0/in_1010 multiplexer_0/in_1011 multiplexer_0/in_1100 multiplexer_0/in_1101
+ multiplexer_0/in_1110 multiplexer_0/in_1111 level_shifter_2/out_b level_shifter_0/out_b
+ avss avdd multiplexer
Xlevel_shifter_0 vtrip[0] level_shifter_0/out level_shifter_0/out_b dvss avss dvdd
+ avdd level_shifter
Xlevel_shifter_1 vtrip[1] level_shifter_1/out level_shifter_1/out_b dvss avss dvdd
+ avdd level_shifter
Xlevel_shifter_2 vtrip[2] level_shifter_2/out level_shifter_2/out_b dvss avss dvdd
+ avdd level_shifter
Xlevel_shifter_3 vtrip[3] level_shifter_3/out level_shifter_3/out_b dvss avss dvdd
+ avdd level_shifter
Xcomp_hyst_0 ovout vbg vin ena ibias dvss dvdd comp_hyst
.ends


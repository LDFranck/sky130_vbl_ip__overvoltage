magic
tech sky130A
magscale 1 2
timestamp 1713226135
<< locali >>
rect 1217 12802 1293 12838
rect 1217 12248 1225 12802
rect 1287 12248 1293 12802
rect 1217 12212 1293 12248
rect 2895 12802 2971 12838
rect 2895 12248 2903 12802
rect 2965 12248 2971 12802
rect 2895 12212 2971 12248
rect 4563 6757 4627 6793
rect 4563 6203 4569 6757
rect 4621 6203 4627 6757
rect 4563 6167 4627 6203
rect 6231 6757 6295 6793
rect 6231 6203 6237 6757
rect 6289 6203 6295 6757
rect 6231 6167 6295 6203
rect 1217 702 1293 738
rect 1217 148 1225 702
rect 1287 148 1293 702
rect 1217 112 1293 148
rect 2895 702 2971 738
rect 2895 148 2903 702
rect 2965 148 2971 702
rect 2895 112 2971 148
<< viali >>
rect 1225 12248 1287 12802
rect 2903 12248 2965 12802
rect 4569 6203 4621 6757
rect 6237 6203 6289 6757
rect 1225 148 1287 702
rect 2903 148 2965 702
<< metal1 >>
rect 1 12910 117 13026
rect 1101 12910 1217 13026
rect 1479 12949 1607 13095
rect 1479 12891 1485 12949
rect 1601 12891 1607 12949
rect 1635 12910 1751 13026
rect 2735 12910 2851 13026
rect 3157 12949 3285 12955
rect 1217 12802 1293 12838
rect 1217 12248 1225 12802
rect 1287 12248 1293 12802
rect 1479 12744 1607 12891
rect 3157 12891 3163 12949
rect 3279 12891 3285 12949
rect 3313 12910 3429 13026
rect 4413 12910 4529 13026
rect 1335 12738 1607 12744
rect 1335 12622 1341 12738
rect 1457 12622 1607 12738
rect 1335 12616 1607 12622
rect 1321 12428 1449 12434
rect 1321 12312 1327 12428
rect 1443 12312 1449 12428
rect 1321 12306 1449 12312
rect 1217 12212 1293 12248
rect 1245 12160 1451 12166
rect 1245 12052 1251 12160
rect 1445 12052 1451 12160
rect 1245 11563 1451 12052
rect 1245 11373 1303 11563
rect 1393 11373 1451 11563
rect 1245 11247 1451 11373
rect 1245 11057 1303 11247
rect 1393 11057 1451 11247
rect 1245 10550 1451 11057
rect 1245 10442 1251 10550
rect 1445 10442 1451 10550
rect 1245 10436 1451 10442
rect 1479 9729 1607 12616
rect 2851 12802 2971 12838
rect 2851 12248 2903 12802
rect 2965 12248 2971 12802
rect 3157 12744 3285 12891
rect 3013 12738 3285 12744
rect 3013 12622 3019 12738
rect 3135 12622 3285 12738
rect 3013 12616 3285 12622
rect 2999 12428 3127 12434
rect 2999 12312 3005 12428
rect 3121 12312 3127 12428
rect 2999 12306 3127 12312
rect 2851 12212 2971 12248
rect 2879 12160 3085 12166
rect 2879 12052 2885 12160
rect 3079 12052 3085 12160
rect 2879 10550 3085 12052
rect 2879 10442 2885 10550
rect 3079 10442 3085 10550
rect 2879 10436 3085 10442
rect 1479 9671 1485 9729
rect 1601 9671 1607 9729
rect 1245 8940 1451 8946
rect 1245 8832 1251 8940
rect 1445 8832 1451 8940
rect 1245 8343 1451 8832
rect 1245 8153 1303 8343
rect 1393 8153 1451 8343
rect 1245 8027 1451 8153
rect 1245 7837 1303 8027
rect 1393 7837 1451 8027
rect 1245 7330 1451 7837
rect 1245 7222 1251 7330
rect 1445 7222 1451 7330
rect 1245 7216 1451 7222
rect 1479 6509 1607 9671
rect 3157 9729 3285 12616
rect 4557 12160 4763 12166
rect 4557 12052 4563 12160
rect 4757 12052 4763 12160
rect 4557 10550 4763 12052
rect 4557 10442 4563 10550
rect 4757 10442 4763 10550
rect 4557 10436 4763 10442
rect 4825 11339 4953 11485
rect 4825 11281 4831 11339
rect 4947 11281 4953 11339
rect 4981 11300 5097 11416
rect 6081 11300 6197 11416
rect 3157 9671 3163 9729
rect 3279 9671 3285 9729
rect 2879 8940 3085 8946
rect 2879 8832 2885 8940
rect 3079 8832 3085 8940
rect 2879 7330 3085 8832
rect 2879 7222 2885 7330
rect 3079 7222 3085 7330
rect 2879 7216 3085 7222
rect 1479 6451 1485 6509
rect 1601 6451 1607 6509
rect 1245 5720 1451 5726
rect 1245 5612 1251 5720
rect 1445 5612 1451 5720
rect 1245 5123 1451 5612
rect 1245 4933 1303 5123
rect 1393 4933 1451 5123
rect 1245 4807 1451 4933
rect 1245 4617 1303 4807
rect 1393 4617 1451 4807
rect 1245 4110 1451 4617
rect 1245 4002 1251 4110
rect 1445 4002 1451 4110
rect 1245 3996 1451 4002
rect 1479 3289 1607 6451
rect 3157 6509 3285 9671
rect 4557 8940 4763 8946
rect 4557 8832 4563 8940
rect 4757 8832 4763 8940
rect 4557 7330 4763 8832
rect 4557 7222 4563 7330
rect 4757 7222 4763 7330
rect 4557 7216 4763 7222
rect 3157 6451 3163 6509
rect 3279 6451 3285 6509
rect 2879 5720 3085 5726
rect 2879 5612 2885 5720
rect 3079 5612 3085 5720
rect 2879 4110 3085 5612
rect 2879 4002 2885 4110
rect 3079 4002 3085 4110
rect 2879 3996 3085 4002
rect 1479 3231 1485 3289
rect 1601 3231 1607 3289
rect 1245 2500 1451 2506
rect 1245 2392 1251 2500
rect 1445 2392 1451 2500
rect 1245 1903 1451 2392
rect 1245 1713 1303 1903
rect 1393 1713 1451 1903
rect 1245 1587 1451 1713
rect 1245 1397 1303 1587
rect 1393 1397 1451 1587
rect 1245 890 1451 1397
rect 1245 782 1251 890
rect 1445 782 1451 890
rect 1245 776 1451 782
rect 1217 702 1293 738
rect 1217 148 1225 702
rect 1287 148 1293 702
rect 1321 638 1449 644
rect 1321 522 1327 638
rect 1443 522 1449 638
rect 1321 516 1449 522
rect 1479 334 1607 3231
rect 3157 3289 3285 6451
rect 4529 6757 4627 6793
rect 4529 6203 4569 6757
rect 4621 6203 4627 6757
rect 4655 6693 4783 6699
rect 4655 6577 4661 6693
rect 4777 6577 4783 6693
rect 4655 6571 4783 6577
rect 4825 6509 4953 11281
rect 6225 10550 6431 10556
rect 6225 10442 6231 10550
rect 6425 10442 6431 10550
rect 4981 8140 5097 9750
rect 6081 8080 6197 9660
rect 6225 7330 6431 10442
rect 6225 7222 6231 7330
rect 6425 7222 6431 7330
rect 6225 7216 6431 7222
rect 6502 8119 6630 8125
rect 6502 8061 6508 8119
rect 6624 8061 6630 8119
rect 6658 8080 6774 8196
rect 7758 8080 7874 8196
rect 4825 6451 4831 6509
rect 4947 6451 4953 6509
rect 4825 6389 4953 6451
rect 4669 6383 4953 6389
rect 4669 6267 4675 6383
rect 4791 6267 4953 6383
rect 4669 6261 4953 6267
rect 4529 6167 4627 6203
rect 4557 5720 4763 5726
rect 4557 5612 4563 5720
rect 4757 5612 4763 5720
rect 4557 4110 4763 5612
rect 4557 4002 4563 4110
rect 4757 4002 4763 4110
rect 4557 3996 4763 4002
rect 3157 3231 3163 3289
rect 3279 3231 3285 3289
rect 2879 2500 3085 2506
rect 2879 2392 2885 2500
rect 3079 2392 3085 2500
rect 2879 890 3085 2392
rect 2879 782 2885 890
rect 3079 782 3085 890
rect 2879 776 3085 782
rect 1335 328 1607 334
rect 1335 212 1341 328
rect 1457 212 1607 328
rect 1335 206 1607 212
rect 1217 112 1293 148
rect 1 -26 117 90
rect 1101 -26 1217 90
rect 1479 69 1607 206
rect 2851 702 2971 738
rect 2851 148 2903 702
rect 2965 148 2971 702
rect 2999 638 3127 644
rect 2999 522 3005 638
rect 3121 522 3127 638
rect 2999 516 3127 522
rect 3157 334 3285 3231
rect 4557 2500 4763 2506
rect 4557 2392 4563 2500
rect 4757 2392 4763 2500
rect 4557 890 4763 2392
rect 4825 1679 4953 6261
rect 6197 6757 6295 6793
rect 6197 6203 6237 6757
rect 6289 6203 6295 6757
rect 6332 6693 6460 6699
rect 6332 6577 6338 6693
rect 6454 6577 6460 6693
rect 6332 6571 6460 6577
rect 6502 6389 6630 8061
rect 6346 6383 6630 6389
rect 6346 6267 6352 6383
rect 6468 6267 6630 6383
rect 6346 6261 6630 6267
rect 6197 6167 6295 6203
rect 6225 5720 6431 5726
rect 6225 5612 6231 5720
rect 6425 5612 6431 5720
rect 4981 3310 5097 4920
rect 6081 2262 6197 4860
rect 6225 2500 6431 5612
rect 6502 4899 6630 6261
rect 7902 7330 8108 7336
rect 7902 7222 7908 7330
rect 8102 7222 8108 7330
rect 7902 5720 8108 7222
rect 7902 5612 7908 5720
rect 8102 5612 8108 5720
rect 7902 5606 8108 5612
rect 6502 4841 6508 4899
rect 6624 4841 6630 4899
rect 6502 4695 6630 4841
rect 6658 4804 6774 4920
rect 7758 4804 7874 4920
rect 6225 2392 6231 2500
rect 6425 2392 6431 2500
rect 6225 2386 6431 2392
rect 4825 1621 4831 1679
rect 4947 1621 4953 1679
rect 4825 1615 4953 1621
rect 4981 1584 5097 1700
rect 6081 1584 6197 1700
rect 4557 782 4563 890
rect 4757 782 4763 890
rect 4557 776 4763 782
rect 3013 328 3285 334
rect 3013 212 3019 328
rect 3135 212 3285 328
rect 3013 206 3285 212
rect 2851 112 2971 148
rect 1479 11 1485 69
rect 1601 11 1607 69
rect 1479 5 1607 11
rect 1635 -26 1751 90
rect 2735 -26 2851 90
rect 3157 69 3285 206
rect 3157 11 3163 69
rect 3279 11 3285 69
rect 3157 -135 3285 11
rect 3313 -26 3429 90
rect 4413 -26 4529 90
<< via1 >>
rect 1485 12891 1601 12949
rect 3163 12891 3279 12949
rect 1341 12622 1457 12738
rect 1327 12312 1443 12428
rect 1251 12052 1445 12160
rect 1303 11373 1393 11563
rect 1303 11057 1393 11247
rect 1251 10442 1445 10550
rect 3019 12622 3135 12738
rect 3005 12312 3121 12428
rect 2885 12052 3079 12160
rect 2885 10442 3079 10550
rect 1485 9671 1601 9729
rect 1251 8832 1445 8940
rect 1303 8153 1393 8343
rect 1303 7837 1393 8027
rect 1251 7222 1445 7330
rect 4563 12052 4757 12160
rect 4563 10442 4757 10550
rect 4831 11281 4947 11339
rect 3163 9671 3279 9729
rect 2885 8832 3079 8940
rect 2885 7222 3079 7330
rect 1485 6451 1601 6509
rect 1251 5612 1445 5720
rect 1303 4933 1393 5123
rect 1303 4617 1393 4807
rect 1251 4002 1445 4110
rect 4563 8832 4757 8940
rect 4563 7222 4757 7330
rect 3163 6451 3279 6509
rect 2885 5612 3079 5720
rect 2885 4002 3079 4110
rect 1485 3231 1601 3289
rect 1251 2392 1445 2500
rect 1303 1713 1393 1903
rect 1303 1397 1393 1587
rect 1251 782 1445 890
rect 1327 522 1443 638
rect 4661 6577 4777 6693
rect 6231 10442 6425 10550
rect 6231 7222 6425 7330
rect 6508 8061 6624 8119
rect 4831 6451 4947 6509
rect 4675 6267 4791 6383
rect 4563 5612 4757 5720
rect 4563 4002 4757 4110
rect 3163 3231 3279 3289
rect 2885 2392 3079 2500
rect 2885 782 3079 890
rect 1341 212 1457 328
rect 3005 522 3121 638
rect 4563 2392 4757 2500
rect 6338 6577 6454 6693
rect 6352 6267 6468 6383
rect 6231 5612 6425 5720
rect 7908 7222 8102 7330
rect 7908 5612 8102 5720
rect 6508 4841 6624 4899
rect 6231 2392 6425 2500
rect 4831 1621 4947 1679
rect 4563 782 4757 890
rect 3019 212 3135 328
rect 1485 11 1601 69
rect 3163 11 3279 69
<< metal2 >>
rect 709 12949 2343 12955
rect 709 12891 1485 12949
rect 1601 12891 2343 12949
rect 709 12885 2343 12891
rect 3157 12949 4021 12955
rect 3157 12891 3163 12949
rect 3279 12891 4021 12949
rect 3157 12885 4021 12891
rect 1335 12738 1463 12744
rect 1335 12622 1341 12738
rect 1457 12622 1463 12738
rect 1335 12616 1463 12622
rect 3013 12738 3141 12744
rect 3013 12622 3019 12738
rect 3135 12622 3141 12738
rect 3013 12616 3141 12622
rect 1307 12439 1463 12448
rect 1307 12301 1316 12439
rect 1454 12301 1463 12439
rect 1307 12292 1463 12301
rect 2985 12439 3141 12448
rect 2985 12301 2994 12439
rect 3132 12301 3141 12439
rect 2985 12292 3141 12301
rect -199 12046 211 12166
rect 1007 12160 1451 12166
rect 1007 12052 1251 12160
rect 1445 12052 1451 12160
rect 1007 12046 1451 12052
rect 1845 12156 2045 12166
rect 1845 12046 2045 12056
rect 2635 12160 3085 12166
rect 2635 12052 2885 12160
rect 3079 12052 3085 12160
rect 2635 12046 3085 12052
rect 3523 12156 3723 12166
rect 3523 12046 3723 12056
rect 4319 12160 4763 12166
rect 4319 12052 4563 12160
rect 4757 12052 4763 12160
rect 4319 12046 4763 12052
rect 1293 11373 1303 11563
rect 1393 11373 1403 11563
rect 709 11339 2343 11345
rect 709 11281 1474 11339
rect 1612 11281 2343 11339
rect 709 11275 2343 11281
rect 3143 11339 4021 11345
rect 3143 11281 3152 11339
rect 3290 11281 4021 11339
rect 3143 11275 4021 11281
rect 4825 11339 5689 11345
rect 4825 11281 4831 11339
rect 4947 11281 5689 11339
rect 4825 11275 5689 11281
rect 1293 11057 1303 11247
rect 1393 11057 1403 11247
rect -199 10436 211 10556
rect 1007 10550 1451 10556
rect 1007 10442 1251 10550
rect 1445 10442 1451 10550
rect 1007 10436 1451 10442
rect 1845 10546 2045 10556
rect 1845 10436 2045 10446
rect 2587 10550 3723 10556
rect 2587 10442 2885 10550
rect 3079 10442 3723 10550
rect 2587 10436 3723 10442
rect 4319 10550 5391 10556
rect 4319 10442 4563 10550
rect 4757 10442 5391 10550
rect 4319 10436 5391 10442
rect 5987 10550 6431 10556
rect 5987 10442 6231 10550
rect 6425 10442 6431 10550
rect 5987 10436 6431 10442
rect 709 9729 2343 9735
rect 709 9671 1485 9729
rect 1601 9671 2343 9729
rect 709 9665 2343 9671
rect 3157 9729 4021 9735
rect 3157 9671 3163 9729
rect 3279 9671 4021 9729
rect 3157 9665 4021 9671
rect 4811 9729 5689 9735
rect 4811 9671 4820 9729
rect 4958 9671 5689 9729
rect 4811 9665 5689 9671
rect -199 8826 211 8946
rect 1007 8940 1451 8946
rect 1007 8832 1251 8940
rect 1445 8832 1451 8940
rect 1007 8826 1451 8832
rect 1845 8936 2045 8946
rect 1845 8826 2045 8836
rect 2641 8940 3085 8946
rect 2641 8832 2885 8940
rect 3079 8832 3085 8940
rect 2641 8826 3085 8832
rect 3523 8936 3723 8946
rect 3523 8826 3723 8836
rect 4319 8940 4763 8946
rect 4319 8832 4563 8940
rect 4757 8832 4763 8940
rect 4319 8826 4763 8832
rect 1293 8153 1303 8343
rect 1393 8153 1403 8343
rect 709 8119 2343 8125
rect 709 8061 1474 8119
rect 1612 8061 2343 8119
rect 709 8055 2343 8061
rect 3143 8119 4021 8125
rect 3143 8061 3152 8119
rect 3290 8061 4021 8119
rect 3143 8055 4021 8061
rect 4811 8119 5689 8125
rect 4811 8061 4820 8119
rect 4958 8061 5689 8119
rect 4811 8055 5689 8061
rect 6502 8119 7366 8125
rect 6502 8061 6508 8119
rect 6624 8061 7366 8119
rect 6502 8055 7366 8061
rect 1293 7837 1303 8027
rect 1393 7837 1403 8027
rect -199 7216 211 7336
rect 1007 7330 1451 7336
rect 1007 7222 1251 7330
rect 1445 7222 1451 7330
rect 1007 7216 1451 7222
rect 1845 7326 2045 7336
rect 1845 7216 2045 7226
rect 2641 7330 3723 7336
rect 2641 7222 2885 7330
rect 3079 7222 3723 7330
rect 2641 7216 3723 7222
rect 4319 7330 5391 7336
rect 4319 7222 4563 7330
rect 4757 7222 5391 7330
rect 4319 7216 5391 7222
rect 5987 7330 7068 7336
rect 5987 7222 6231 7330
rect 6425 7222 7068 7330
rect 5987 7216 7068 7222
rect 7664 7330 8108 7336
rect 7664 7222 7908 7330
rect 8102 7222 8108 7330
rect 7664 7216 8108 7222
rect 4641 6704 4797 6713
rect 4641 6566 4650 6704
rect 4788 6566 4797 6704
rect 4641 6557 4797 6566
rect 6318 6704 6474 6713
rect 6318 6566 6327 6704
rect 6465 6566 6474 6704
rect 6318 6557 6474 6566
rect 709 6509 2343 6515
rect 709 6451 1485 6509
rect 1601 6451 2343 6509
rect 709 6445 2343 6451
rect 3157 6509 4021 6515
rect 3157 6451 3163 6509
rect 3279 6451 4021 6509
rect 3157 6445 4021 6451
rect 4825 6509 5689 6515
rect 4825 6451 4831 6509
rect 4947 6451 5689 6509
rect 4825 6445 5689 6451
rect 6488 6509 7366 6515
rect 6488 6451 6497 6509
rect 6635 6451 7366 6509
rect 6488 6445 7366 6451
rect 4669 6383 4797 6389
rect 4669 6267 4675 6383
rect 4791 6267 4797 6383
rect 4669 6261 4797 6267
rect 6346 6383 6474 6389
rect 6346 6267 6352 6383
rect 6468 6267 6474 6383
rect 6346 6261 6474 6267
rect -199 5606 211 5726
rect 1007 5720 1451 5726
rect 1007 5612 1251 5720
rect 1445 5612 1451 5720
rect 1007 5606 1451 5612
rect 1845 5716 2045 5726
rect 1845 5606 2045 5616
rect 2641 5720 3085 5726
rect 2641 5612 2885 5720
rect 3079 5612 3085 5720
rect 2641 5606 3085 5612
rect 3523 5716 3723 5726
rect 3523 5606 3723 5616
rect 4319 5720 5391 5726
rect 4319 5612 4563 5720
rect 4757 5612 5391 5720
rect 4319 5606 5391 5612
rect 5987 5720 7068 5726
rect 5987 5612 6231 5720
rect 6425 5612 7068 5720
rect 5987 5606 7068 5612
rect 7664 5720 8108 5726
rect 7664 5612 7908 5720
rect 8102 5612 8108 5720
rect 7664 5606 8108 5612
rect 1293 4933 1303 5123
rect 1393 4933 1403 5123
rect 709 4899 2343 4905
rect 709 4841 1474 4899
rect 1612 4841 2343 4899
rect 709 4835 2343 4841
rect 3143 4899 4021 4905
rect 3143 4841 3152 4899
rect 3290 4841 4021 4899
rect 3143 4835 4021 4841
rect 4811 4899 5689 4905
rect 4811 4841 4820 4899
rect 4958 4841 5689 4899
rect 4811 4835 5689 4841
rect 6502 4899 7366 4905
rect 6502 4841 6508 4899
rect 6624 4841 7366 4899
rect 6502 4835 7366 4841
rect 1293 4617 1303 4807
rect 1393 4617 1403 4807
rect -199 3996 211 4116
rect 1007 4110 1451 4116
rect 1007 4002 1251 4110
rect 1445 4002 1451 4110
rect 1007 3996 1451 4002
rect 1845 4106 2045 4116
rect 1845 3996 2045 4006
rect 2641 4110 3723 4116
rect 2641 4002 2885 4110
rect 3079 4002 3723 4110
rect 2641 3996 3723 4002
rect 4319 4110 4763 4116
rect 4319 4002 4563 4110
rect 4757 4002 4763 4110
rect 4319 3996 4763 4002
rect 709 3289 2343 3295
rect 709 3231 1485 3289
rect 1601 3231 2343 3289
rect 709 3225 2343 3231
rect 3157 3289 4021 3295
rect 3157 3231 3163 3289
rect 3279 3231 4021 3289
rect 3157 3225 4021 3231
rect 4811 3289 5689 3295
rect 4811 3231 4820 3289
rect 4958 3231 5689 3289
rect 4811 3225 5689 3231
rect -199 2386 211 2506
rect 1007 2500 1451 2506
rect 1007 2392 1251 2500
rect 1445 2392 1451 2500
rect 1007 2386 1451 2392
rect 1845 2496 2045 2506
rect 1845 2386 2045 2396
rect 2641 2500 3085 2506
rect 2641 2392 2885 2500
rect 3079 2392 3085 2500
rect 2641 2386 3085 2392
rect 3523 2496 3723 2506
rect 3523 2386 3723 2396
rect 4319 2500 5391 2506
rect 4319 2392 4563 2500
rect 4757 2392 5391 2500
rect 4319 2386 5391 2392
rect 5987 2500 6431 2506
rect 5987 2392 6231 2500
rect 6425 2392 6431 2500
rect 5987 2386 6431 2392
rect 1293 1713 1303 1903
rect 1393 1713 1403 1903
rect 709 1679 2343 1685
rect 709 1621 1474 1679
rect 1612 1621 2343 1679
rect 709 1615 2343 1621
rect 3143 1679 4021 1685
rect 3143 1621 3152 1679
rect 3290 1621 4021 1679
rect 3143 1615 4021 1621
rect 4825 1679 5689 1685
rect 4825 1621 4831 1679
rect 4947 1621 5689 1679
rect 4825 1615 5689 1621
rect 1293 1397 1303 1587
rect 1393 1397 1403 1587
rect -199 776 211 896
rect 1007 890 1451 896
rect 1007 782 1251 890
rect 1445 782 1451 890
rect 1007 776 1451 782
rect 1845 886 2045 896
rect 1845 776 2045 786
rect 2641 890 3723 896
rect 2641 782 2885 890
rect 3079 782 3723 890
rect 2641 776 3723 782
rect 4319 890 4763 896
rect 4319 782 4563 890
rect 4757 782 4763 890
rect 4319 776 4763 782
rect 1307 649 1463 658
rect 1307 511 1316 649
rect 1454 511 1463 649
rect 1307 502 1463 511
rect 2985 649 3141 658
rect 2985 511 2994 649
rect 3132 511 3141 649
rect 2985 502 3141 511
rect 1335 328 1463 334
rect 1335 212 1341 328
rect 1457 212 1463 328
rect 1335 206 1463 212
rect 3013 328 3141 334
rect 3013 212 3019 328
rect 3135 212 3141 328
rect 3013 206 3141 212
rect 709 69 2343 75
rect 709 11 1485 69
rect 1601 11 2343 69
rect 709 5 2343 11
rect 3157 69 4021 75
rect 3157 11 3163 69
rect 3279 11 4021 69
rect 3157 5 4021 11
<< via2 >>
rect 1316 12428 1454 12439
rect 1316 12312 1327 12428
rect 1327 12312 1443 12428
rect 1443 12312 1454 12428
rect 1316 12301 1454 12312
rect 2994 12428 3132 12439
rect 2994 12312 3005 12428
rect 3005 12312 3121 12428
rect 3121 12312 3132 12428
rect 2994 12301 3132 12312
rect 1845 12056 2045 12156
rect 3523 12056 3723 12156
rect 1303 11373 1393 11563
rect 1474 11281 1612 11339
rect 3152 11281 3290 11339
rect 1303 11057 1393 11247
rect 1845 10446 2045 10546
rect 4820 9671 4958 9729
rect 1845 8836 2045 8936
rect 3523 8836 3723 8936
rect 1303 8153 1393 8343
rect 1474 8061 1612 8119
rect 3152 8061 3290 8119
rect 4820 8061 4958 8119
rect 1303 7837 1393 8027
rect 1845 7226 2045 7326
rect 4650 6693 4788 6704
rect 4650 6577 4661 6693
rect 4661 6577 4777 6693
rect 4777 6577 4788 6693
rect 4650 6566 4788 6577
rect 6327 6693 6465 6704
rect 6327 6577 6338 6693
rect 6338 6577 6454 6693
rect 6454 6577 6465 6693
rect 6327 6566 6465 6577
rect 6497 6451 6635 6509
rect 1845 5616 2045 5716
rect 3523 5616 3723 5716
rect 1303 4933 1393 5123
rect 1474 4841 1612 4899
rect 3152 4841 3290 4899
rect 4820 4841 4958 4899
rect 1303 4617 1393 4807
rect 1845 4006 2045 4106
rect 4820 3231 4958 3289
rect 1845 2396 2045 2496
rect 3523 2396 3723 2496
rect 1303 1713 1393 1903
rect 1474 1621 1612 1679
rect 3152 1621 3290 1679
rect 1303 1397 1393 1587
rect 1845 786 2045 886
rect 1316 638 1454 649
rect 1316 522 1327 638
rect 1327 522 1443 638
rect 1443 522 1454 638
rect 1316 511 1454 522
rect 2994 638 3132 649
rect 2994 522 3005 638
rect 3005 522 3121 638
rect 3121 522 3132 638
rect 2994 511 3132 522
<< metal3 >>
rect 1469 12448 1617 13025
rect 3147 12448 3295 12955
rect 1307 12439 1617 12448
rect 1307 12301 1316 12439
rect 1454 12301 1617 12439
rect 1307 12292 1617 12301
rect 2985 12439 3295 12448
rect 2985 12301 2994 12439
rect 3132 12301 3295 12439
rect 2985 12292 3295 12301
rect 1298 11563 1398 11573
rect 1298 11373 1303 11563
rect 1393 11373 1398 11563
rect 1298 11363 1398 11373
rect 1469 11339 1617 12292
rect 1835 12156 2055 12161
rect 1835 12056 1845 12156
rect 2045 12056 2055 12156
rect 1835 12051 2055 12056
rect 2877 12060 2887 12150
rect 3077 12060 3087 12150
rect 1469 11281 1474 11339
rect 1612 11281 1617 11339
rect 1298 11247 1398 11257
rect 1298 11057 1303 11247
rect 1393 11057 1398 11247
rect 1298 11047 1398 11057
rect 1298 8343 1398 8353
rect 1298 8153 1303 8343
rect 1393 8153 1398 8343
rect 1298 8143 1398 8153
rect 1469 8119 1617 11281
rect 2877 11355 3087 12060
rect 2877 11265 2887 11355
rect 3077 11265 3087 11355
rect 3147 11339 3295 12292
rect 3513 12156 3733 12161
rect 3513 12056 3523 12156
rect 3723 12056 3733 12156
rect 3513 12051 3733 12056
rect 4816 11345 4963 11415
rect 3147 11281 3152 11339
rect 3290 11281 3295 11339
rect 1835 10546 2055 10551
rect 1835 10446 1845 10546
rect 2045 10446 2055 10546
rect 1835 10441 2055 10446
rect 1835 8936 2055 8941
rect 1835 8836 1845 8936
rect 2045 8836 2055 8936
rect 1835 8831 2055 8836
rect 2877 8840 2887 8930
rect 3077 8840 3087 8930
rect 1469 8061 1474 8119
rect 1612 8061 1617 8119
rect 1298 8027 1398 8037
rect 1298 7837 1303 8027
rect 1393 7837 1398 8027
rect 1298 7827 1398 7837
rect 1298 5123 1398 5133
rect 1298 4933 1303 5123
rect 1393 4933 1398 5123
rect 1298 4923 1398 4933
rect 1469 4899 1617 8061
rect 2877 8135 3087 8840
rect 2877 8045 2887 8135
rect 3077 8045 3087 8135
rect 3147 8119 3295 11281
rect 4815 9729 4963 11345
rect 4815 9671 4820 9729
rect 4958 9671 4963 9729
rect 3513 8936 3733 8941
rect 3513 8836 3523 8936
rect 3723 8836 3733 8936
rect 3513 8831 3733 8836
rect 3147 8061 3152 8119
rect 3290 8061 3295 8119
rect 1835 7326 2055 7331
rect 1835 7226 1845 7326
rect 2045 7226 2055 7326
rect 1835 7221 2055 7226
rect 1835 5716 2055 5721
rect 1835 5616 1845 5716
rect 2045 5616 2055 5716
rect 1835 5611 2055 5616
rect 2877 5620 2887 5710
rect 3077 5620 3087 5710
rect 1469 4841 1474 4899
rect 1612 4841 1617 4899
rect 1298 4807 1398 4817
rect 1298 4617 1303 4807
rect 1393 4617 1398 4807
rect 1298 4607 1398 4617
rect 1298 1903 1398 1913
rect 1298 1713 1303 1903
rect 1393 1713 1398 1903
rect 1298 1703 1398 1713
rect 1469 1679 1617 4841
rect 2877 4915 3087 5620
rect 2877 4825 2887 4915
rect 3077 4825 3087 4915
rect 3147 4899 3295 8061
rect 4815 8119 4963 9671
rect 4815 8061 4820 8119
rect 4958 8061 4963 8119
rect 4815 6713 4963 8061
rect 6492 6713 6640 8125
rect 4641 6704 4963 6713
rect 4641 6566 4650 6704
rect 4788 6566 4963 6704
rect 4641 6557 4963 6566
rect 6318 6704 6640 6713
rect 6318 6566 6327 6704
rect 6465 6566 6640 6704
rect 6318 6557 6640 6566
rect 3513 5716 3733 5721
rect 3513 5616 3523 5716
rect 3723 5616 3733 5716
rect 3513 5611 3733 5616
rect 3147 4841 3152 4899
rect 3290 4841 3295 4899
rect 1835 4106 2055 4111
rect 1835 4006 1845 4106
rect 2045 4006 2055 4106
rect 1835 4001 2055 4006
rect 1835 2496 2055 2501
rect 1835 2396 1845 2496
rect 2045 2396 2055 2496
rect 1835 2391 2055 2396
rect 2877 2400 2887 2490
rect 3077 2400 3087 2490
rect 1469 1621 1474 1679
rect 1612 1621 1617 1679
rect 1298 1587 1398 1597
rect 1298 1397 1303 1587
rect 1393 1397 1398 1587
rect 1298 1387 1398 1397
rect 1469 658 1617 1621
rect 2877 1695 3087 2400
rect 2877 1605 2887 1695
rect 3077 1605 3087 1695
rect 3147 1679 3295 4841
rect 4815 4899 4963 6557
rect 4815 4841 4820 4899
rect 4958 4841 4963 4899
rect 4815 3289 4963 4841
rect 6492 6509 6640 6557
rect 6492 6451 6497 6509
rect 6635 6451 6640 6509
rect 6492 4765 6640 6451
rect 4815 3231 4820 3289
rect 4958 3231 4963 3289
rect 3513 2496 3733 2501
rect 3513 2396 3523 2496
rect 3723 2396 3733 2496
rect 3513 2391 3733 2396
rect 3147 1621 3152 1679
rect 3290 1621 3295 1679
rect 1835 886 2055 891
rect 1835 786 1845 886
rect 2045 786 2055 886
rect 1835 781 2055 786
rect 3147 658 3295 1621
rect 4815 1615 4963 3231
rect 1307 649 1617 658
rect 1307 511 1316 649
rect 1454 511 1617 649
rect 1307 502 1617 511
rect 2985 649 3295 658
rect 2985 511 2994 649
rect 3132 511 3295 649
rect 2985 502 3295 511
rect 1469 5 1617 502
rect 3147 -65 3295 502
<< via3 >>
rect 1303 11373 1393 11563
rect 1845 12056 2045 12156
rect 2887 12060 3077 12150
rect 1303 11057 1393 11247
rect 1303 8153 1393 8343
rect 2887 11265 3077 11355
rect 3523 12056 3723 12156
rect 1845 10446 2045 10546
rect 1845 8836 2045 8936
rect 2887 8840 3077 8930
rect 1303 7837 1393 8027
rect 1303 4933 1393 5123
rect 2887 8045 3077 8135
rect 3523 8836 3723 8936
rect 1845 7226 2045 7326
rect 1845 5616 2045 5716
rect 2887 5620 3077 5710
rect 1303 4617 1393 4807
rect 1303 1713 1393 1903
rect 2887 4825 3077 4915
rect 3523 5616 3723 5716
rect 1845 4006 2045 4106
rect 1845 2396 2045 2496
rect 2887 2400 3077 2490
rect 1303 1397 1393 1587
rect 2887 1605 3077 1695
rect 3523 2396 3723 2496
rect 1845 786 2045 886
<< metal4 >>
rect -99 12156 2046 12157
rect -99 12056 1845 12156
rect 2045 12056 2046 12156
rect -99 12055 2046 12056
rect 2882 12156 3724 12157
rect 2882 12150 3523 12156
rect 2882 12060 2887 12150
rect 3077 12060 3523 12150
rect 2882 12056 3523 12060
rect 3723 12056 3724 12156
rect 2882 12055 3724 12056
rect 1298 11563 1398 11568
rect 1298 11373 1303 11563
rect 1393 11373 1398 11563
rect 1298 11360 1398 11373
rect 1298 11355 3082 11360
rect 1298 11265 2887 11355
rect 3077 11265 3082 11355
rect 1298 11260 3082 11265
rect 1298 11247 1398 11260
rect 1298 11057 1303 11247
rect 1393 11057 1398 11247
rect 1298 11052 1398 11057
rect -99 10546 2046 10547
rect -99 10446 1845 10546
rect 2045 10446 2046 10546
rect -99 10445 2046 10446
rect -99 8936 2046 8937
rect -99 8836 1845 8936
rect 2045 8836 2046 8936
rect -99 8835 2046 8836
rect 2882 8936 3724 8937
rect 2882 8930 3523 8936
rect 2882 8840 2887 8930
rect 3077 8840 3523 8930
rect 2882 8836 3523 8840
rect 3723 8836 3724 8936
rect 2882 8835 3724 8836
rect 1298 8343 1398 8348
rect 1298 8153 1303 8343
rect 1393 8153 1398 8343
rect 1298 8140 1398 8153
rect 1298 8135 3082 8140
rect 1298 8045 2887 8135
rect 3077 8045 3082 8135
rect 1298 8040 3082 8045
rect 1298 8027 1398 8040
rect 1298 7837 1303 8027
rect 1393 7837 1398 8027
rect 1298 7832 1398 7837
rect -99 7326 2046 7327
rect -99 7226 1845 7326
rect 2045 7226 2046 7326
rect -99 7225 2046 7226
rect -99 5716 2046 5717
rect -99 5616 1845 5716
rect 2045 5616 2046 5716
rect -99 5615 2046 5616
rect 2882 5716 3724 5717
rect 2882 5710 3523 5716
rect 2882 5620 2887 5710
rect 3077 5620 3523 5710
rect 2882 5616 3523 5620
rect 3723 5616 3724 5716
rect 2882 5615 3724 5616
rect 1298 5123 1398 5128
rect 1298 4933 1303 5123
rect 1393 4933 1398 5123
rect 1298 4920 1398 4933
rect 1298 4915 3082 4920
rect 1298 4825 2887 4915
rect 3077 4825 3082 4915
rect 1298 4820 3082 4825
rect 1298 4807 1398 4820
rect 1298 4617 1303 4807
rect 1393 4617 1398 4807
rect 1298 4612 1398 4617
rect -99 4106 2046 4107
rect -99 4006 1845 4106
rect 2045 4006 2046 4106
rect -99 4005 2046 4006
rect -99 2496 2046 2497
rect -99 2396 1845 2496
rect 2045 2396 2046 2496
rect -99 2395 2046 2396
rect 2882 2496 3724 2497
rect 2882 2490 3523 2496
rect 2882 2400 2887 2490
rect 3077 2400 3523 2490
rect 2882 2396 3523 2400
rect 3723 2396 3724 2496
rect 2882 2395 3724 2396
rect 1298 1903 1398 1908
rect 1298 1713 1303 1903
rect 1393 1713 1398 1903
rect 1298 1700 1398 1713
rect 1298 1695 3082 1700
rect 1298 1605 2887 1695
rect 3077 1605 3082 1695
rect 1298 1600 3082 1605
rect 1298 1587 1398 1600
rect 1298 1397 1303 1587
rect 1393 1397 1398 1587
rect 1298 1392 1398 1397
rect -99 886 2046 887
rect -99 786 1845 886
rect 2045 786 2046 886
rect -99 785 2046 786
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_0
timestamp 1713221383
transform 1 0 1406 0 1 12680
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_1
timestamp 1713221383
transform 1 0 1406 0 1 12370
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_2
timestamp 1713221383
transform 1 0 1406 0 -1 580
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_3
timestamp 1713221383
transform 1 0 1406 0 -1 270
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_4
timestamp 1713221383
transform 1 0 3084 0 -1 270
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_5
timestamp 1713221383
transform 1 0 3084 0 -1 580
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_6
timestamp 1713221383
transform 1 0 3084 0 1 12370
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_7
timestamp 1713221383
transform 1 0 3084 0 1 12680
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_8
timestamp 1713221383
transform 1 0 4740 0 -1 6635
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_9
timestamp 1713221383
transform 1 0 4740 0 -1 6325
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_10
timestamp 1713221383
transform 1 0 6417 0 -1 6635
box -183 -208 183 208
use sky130_fd_pr__diode_pw2nd_05v5_F6RBXN  sky130_fd_pr__diode_pw2nd_05v5_F6RBXN_11
timestamp 1713221383
transform 1 0 6417 0 -1 6325
box -183 -208 183 208
use trans_gate_m  trans_gate_m_0
timestamp 1713221383
transform 1 0 1780 0 1 11415
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_1
timestamp 1713221383
transform 1 0 1780 0 1 9805
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_2
timestamp 1713221383
transform 1 0 1780 0 1 8195
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_3
timestamp 1713221383
transform 1 0 1780 0 1 6585
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_4
timestamp 1713221383
transform 1 0 1780 0 1 3365
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_5
timestamp 1713221383
transform 1 0 1780 0 1 4975
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_6
timestamp 1713221383
transform 1 0 1780 0 1 1755
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_7
timestamp 1713221383
transform 1 0 1780 0 1 145
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_8
timestamp 1713221383
transform 1 0 146 0 1 145
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_9
timestamp 1713221383
transform 1 0 146 0 1 1755
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_10
timestamp 1713221383
transform 1 0 146 0 1 4975
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_11
timestamp 1713221383
transform 1 0 146 0 1 3365
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_12
timestamp 1713221383
transform 1 0 146 0 1 6585
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_13
timestamp 1713221383
transform 1 0 146 0 1 8195
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_14
timestamp 1713221383
transform 1 0 146 0 1 9805
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_15
timestamp 1713221383
transform 1 0 146 0 1 11415
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_18
timestamp 1713221383
transform 1 0 3458 0 1 1755
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_19
timestamp 1713221383
transform 1 0 3458 0 1 145
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_20
timestamp 1713221383
transform 1 0 5126 0 1 9805
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_21
timestamp 1713221383
transform 1 0 3458 0 1 3365
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_23
timestamp 1713221383
transform 1 0 3458 0 1 4975
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_25
timestamp 1713221383
transform 1 0 3458 0 1 6585
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_27
timestamp 1713221383
transform 1 0 3458 0 1 8195
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_28
timestamp 1713221383
transform 1 0 5126 0 1 6585
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_29
timestamp 1713221383
transform 1 0 3458 0 1 9805
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_31
timestamp 1713221383
transform 1 0 3458 0 1 11415
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_32
timestamp 1713221383
transform 1 0 5126 0 1 4975
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_33
timestamp 1713221383
transform 1 0 6803 0 1 6585
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_34
timestamp 1713221383
transform 1 0 6803 0 1 4975
box -145 -145 1071 1555
use trans_gate_m  trans_gate_m_37
timestamp 1713221383
transform 1 0 5126 0 1 1755
box -145 -145 1071 1555
<< labels >>
flabel metal2 -199 2396 -99 2496 7 FreeSans 800 0 0 0 in_1100
port 24 w
flabel metal2 -199 786 -99 886 7 FreeSans 800 0 0 0 in_1101
port 25 w
flabel metal2 -199 4006 -99 4106 7 FreeSans 800 0 0 0 in_1001
port 21 w
flabel metal2 -199 5616 -99 5716 7 FreeSans 800 0 0 0 in_1000
port 20 w
flabel metal2 -199 7226 -99 7326 7 FreeSans 800 0 0 0 in_0101
port 6 w
flabel metal2 -199 8836 -99 8936 7 FreeSans 800 0 0 0 in_0100
port 5 w
flabel metal2 -199 10446 -99 10546 7 FreeSans 800 0 0 0 in_0001
port 2 w
flabel metal2 -199 12056 -99 12156 7 FreeSans 800 0 0 0 in_0000
port 1 w
flabel metal4 -99 786 1 886 3 FreeSans 800 0 0 0 in_1111
port 27 e
flabel metal4 -99 2396 1 2496 3 FreeSans 800 0 0 0 in_1110
port 26 e
flabel metal4 -99 4006 1 4106 3 FreeSans 800 0 0 0 in_1011
port 23 e
flabel metal4 -99 5616 1 5716 3 FreeSans 800 0 0 0 in_1010
port 22 e
flabel metal4 -99 7226 1 7326 3 FreeSans 800 0 0 0 in_0111
port 10 e
flabel metal4 -99 8836 1 8936 3 FreeSans 800 0 0 0 in_0110
port 7 e
flabel metal4 -99 10446 1 10546 3 FreeSans 800 0 0 0 in_0011
port 4 e
flabel metal4 -99 12056 1 12156 3 FreeSans 800 0 0 0 in_0010
port 3 e
flabel metal1 1508 13025 1578 13095 0 FreeSans 800 0 0 0 vtrip_0
port 18 nsew
flabel metal3 1508 12955 1578 13025 0 FreeSans 800 0 0 0 vtrip_0_b
port 19 nsew
flabel metal1 1131 12970 1187 13026 0 FreeSans 800 0 0 0 vss
port 9 nsew
flabel metal1 31 12970 87 13026 0 FreeSans 800 0 0 0 avdd
port 8 nsew
flabel metal1 1665 12970 1721 13026 0 FreeSans 800 0 0 0 avdd
flabel metal1 2765 12970 2821 13026 0 FreeSans 800 0 0 0 vss
flabel metal1 3343 12970 3399 13026 0 FreeSans 800 0 0 0 avdd
flabel metal1 4443 12970 4499 13026 0 FreeSans 800 0 0 0 vss
flabel metal3 3186 -65 3256 5 0 FreeSans 800 0 0 0 vtrip_1_b
port 17 nsew
flabel metal1 3186 -135 3256 -65 0 FreeSans 800 0 0 0 vtrip_1
port 15 nsew
flabel metal1 5011 11360 5067 11416 0 FreeSans 800 0 0 0 avdd
flabel metal1 6111 11360 6167 11416 0 FreeSans 800 0 0 0 vss
flabel metal1 4854 11415 4924 11485 0 FreeSans 800 0 0 0 vtrip_2
port 13 nsew
flabel metal3 4854 11345 4924 11415 0 FreeSans 800 0 0 0 vtrip_2_b
port 14 nsew
flabel metal1 6531 4695 6601 4765 0 FreeSans 800 0 0 0 vtrip_3
port 11 nsew
flabel metal3 6531 4765 6601 4835 0 FreeSans 800 0 0 0 vtrip_3_b
port 12 nsew
flabel metal1 6688 8140 6744 8196 0 FreeSans 800 0 0 0 avdd
flabel metal1 7788 8140 7844 8196 0 FreeSans 800 0 0 0 vss
flabel metal1 8008 6430 8108 6530 0 FreeSans 800 0 0 0 out
port 16 nsew
<< end >>

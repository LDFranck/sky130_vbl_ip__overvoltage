** sch_path: /home/vblabs/sky130_vbl_ip__overvoltage/blocks/comp_hyst/xschem/comp_hyst.sch
.subckt comp_hyst dvdd out vref vin ena ibias vss
*.PININFO dvdd:B vref:I vin:I out:O ibias:I ena:I vss:B
XM5[0] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM5[1] net3 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM3[0] net4 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM3[1] net4 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM7 net2 net4 dvdd dvdd sky130_fd_pr__pfet_01v8 L=8 W=1 nf=1 m=1
XM4[0] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM4[1] net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM11 net5 net5 vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM12 net1 net5 vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 m=1
XM9 out net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 m=1
XM10 out net2 vss vss sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 m=1
XM17 out ena_b vss vss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM1[0] net4 vref net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM1[1] net4 vref net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM2[0] net3 vin net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM2[1] net3 vin net1 vss sky130_fd_pr__nfet_g5v0d10v5 L=8 W=1.3 nf=1 m=1
XM13 net5 ena_b vss vss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM6[0] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM6[1] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM6[2] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM6[3] net4 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=16 W=1 nf=1 m=1
XM8 net2 net2 vss vss sky130_fd_pr__nfet_01v8 L=8 W=1 nf=1 m=1
XM16 net3 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM15 net4 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM14 net2 ena_b vss vss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
XM18 ena_b ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 m=1
XM19 ena_b ena vss vss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 m=1
x1 ibias ena_b ena dvdd vss net5 trans_gate
.ends

* expanding   symbol:  trans_gate.sym # of pins=6
** sym_path: /home/vblabs/sky130_vbl_ip__overvoltage/blocks/comp_hyst/xschem/trans_gate.sym
** sch_path: /home/vblabs/sky130_vbl_ip__overvoltage/blocks/comp_hyst/xschem/trans_gate.sch
.subckt trans_gate in ena_b ena avdd vss out
*.PININFO avdd:B vss:B ena:I ena_b:I in:I out:I
XM1 in ena out vss sky130_fd_pr__nfet_g5v0d10v5 L=5 W=1 nf=1 m=1
XM2 in ena_b out avdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=6 nf=1 m=1
.ends

.end

magic
tech sky130A
timestamp 1713221383
<< pwell >>
rect -514 -194 514 194
<< mvnmos >>
rect -400 -65 400 65
<< mvndiff >>
rect -429 59 -400 65
rect -429 -59 -423 59
rect -406 -59 -400 59
rect -429 -65 -400 -59
rect 400 59 429 65
rect 400 -59 406 59
rect 423 -59 429 59
rect 400 -65 429 -59
<< mvndiffc >>
rect -423 -59 -406 59
rect 406 -59 423 59
<< mvpsubdiff >>
rect -496 170 496 176
rect -496 153 -442 170
rect 442 153 496 170
rect -496 147 496 153
rect -496 122 -467 147
rect -496 -122 -490 122
rect -473 -122 -467 122
rect 467 122 496 147
rect -496 -147 -467 -122
rect 467 -122 473 122
rect 490 -122 496 122
rect 467 -147 496 -122
rect -496 -153 496 -147
rect -496 -170 -442 -153
rect 442 -170 496 -153
rect -496 -176 496 -170
<< mvpsubdiffcont >>
rect -442 153 442 170
rect -490 -122 -473 122
rect 473 -122 490 122
rect -442 -170 442 -153
<< poly >>
rect -400 101 400 109
rect -400 84 -392 101
rect 392 84 400 101
rect -400 65 400 84
rect -400 -84 400 -65
rect -400 -101 -392 -84
rect 392 -101 400 -84
rect -400 -109 400 -101
<< polycont >>
rect -392 84 392 101
rect -392 -101 392 -84
<< locali >>
rect -490 153 -442 170
rect 442 153 490 170
rect -490 122 -473 153
rect 473 122 490 153
rect -400 84 -392 101
rect 392 84 400 101
rect -423 59 -406 67
rect -423 -67 -406 -59
rect 406 59 423 67
rect 406 -67 423 -59
rect -400 -101 -392 -84
rect 392 -101 400 -84
rect -490 -153 -473 -122
rect 473 -153 490 -122
rect -490 -170 -442 -153
rect 442 -170 490 -153
<< viali >>
rect -392 84 392 101
rect -423 -59 -406 59
rect 406 -59 423 59
rect -392 -101 392 -84
<< metal1 >>
rect -398 101 398 104
rect -398 84 -392 101
rect 392 84 398 101
rect -398 81 398 84
rect -426 59 -403 65
rect -426 -59 -423 59
rect -406 -59 -403 59
rect -426 -65 -403 -59
rect 403 59 426 65
rect 403 -59 406 59
rect 423 -59 426 59
rect 403 -65 426 -59
rect -398 -84 398 -81
rect -398 -101 -392 -84
rect 392 -101 398 -84
rect -398 -104 398 -101
<< properties >>
string FIXED_BBOX -481 -161 481 161
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1.3 l 8.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

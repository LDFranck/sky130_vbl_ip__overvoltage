magic
tech sky130A
magscale 1 2
timestamp 1712255915
<< nwell >>
rect 25583 1972 25585 1974
rect 25645 1972 25647 1974
rect 25326 1662 25402 1865
rect 15090 -22 15108 -7
rect 15090 -26 15151 -22
rect 15090 -54 15108 -26
rect 14668 -1650 14880 -1603
<< poly >>
rect 25645 1972 25647 1974
<< metal1 >>
rect 21308 2762 25871 2808
rect 21308 2480 21354 2762
rect 21566 2480 21612 2762
rect 21794 2480 21841 2762
rect 23452 2480 23499 2762
rect 23680 2480 23727 2762
rect 25339 2480 25386 2762
rect 25566 2480 25612 2762
rect 25825 2480 25871 2762
rect 21308 2434 25871 2480
rect 21308 2276 21354 2434
rect 21566 2276 21612 2434
rect 21308 2230 21612 2276
rect 21308 1948 21354 2230
rect 21566 1948 21612 2230
rect 21778 1989 21788 2189
rect 21840 1989 21850 2189
rect 22418 1948 22815 2277
rect 23504 2189 23673 2434
rect 23453 1989 23726 2189
rect 24340 1948 24737 2277
rect 25566 2276 25612 2434
rect 25825 2276 25871 2434
rect 25566 2230 25871 2276
rect 25328 1989 25338 2189
rect 25390 1989 25400 2189
rect 25566 1948 25612 2230
rect 25825 1948 25871 2230
rect 21308 1902 21612 1948
rect 21308 1744 21354 1902
rect 21566 1744 21612 1902
rect 21308 1698 21612 1744
rect 21850 1698 25327 1948
rect 25566 1902 25871 1948
rect 25566 1744 25612 1902
rect 25825 1744 25871 1902
rect 25566 1698 25871 1744
rect 21308 1416 21354 1698
rect 21566 1416 21612 1698
rect 21778 1458 21788 1657
rect 21840 1458 21850 1657
rect 21308 1370 21612 1416
rect 21308 1212 21354 1370
rect 21566 1212 21612 1370
rect 22418 1369 22815 1698
rect 23451 1457 23726 1657
rect 23499 1212 23668 1457
rect 24339 1370 24736 1698
rect 25328 1456 25338 1657
rect 25390 1456 25400 1657
rect 25566 1416 25612 1698
rect 25825 1416 25871 1698
rect 25566 1370 25871 1416
rect 25566 1212 25612 1370
rect 25825 1212 25871 1370
rect 21308 1166 25871 1212
rect 21308 884 21354 1166
rect 21566 884 21612 1166
rect 21794 884 21841 1166
rect 23452 884 23499 1166
rect 23680 884 23727 1166
rect 25338 884 25385 1166
rect 25566 884 25612 1166
rect 25825 884 25871 1166
rect 21308 838 25871 884
rect 14622 273 25870 320
rect 14622 -7 14668 273
rect 14880 -7 14926 273
rect 15108 -7 15154 273
rect 25566 -7 25612 273
rect 25824 -7 25870 273
rect 14622 -54 25870 -7
rect 14622 -55 14926 -54
rect 14622 -211 14668 -55
rect 14880 -211 14926 -55
rect 14622 -258 14926 -211
rect 14622 -539 14668 -258
rect 14880 -299 14926 -258
rect 14880 -499 15154 -299
rect 14880 -539 14926 -499
rect 14622 -586 14926 -539
rect 16580 -540 16976 -211
rect 18356 -499 18366 -299
rect 18418 -499 18428 -299
rect 18538 -500 18622 -54
rect 20120 -540 20516 -210
rect 21842 -499 21852 -299
rect 21904 -499 21914 -299
rect 22064 -499 22074 -299
rect 22126 -499 22136 -299
rect 23640 -540 24036 -210
rect 25566 -211 25612 -54
rect 25824 -211 25870 -54
rect 25566 -258 25870 -211
rect 25566 -299 25612 -258
rect 25338 -499 25612 -299
rect 25566 -539 25612 -499
rect 25824 -539 25870 -258
rect 14622 -743 14668 -586
rect 14880 -743 14926 -586
rect 14622 -790 14926 -743
rect 15164 -790 25328 -540
rect 25566 -586 25870 -539
rect 25566 -743 25612 -586
rect 25824 -743 25870 -586
rect 25566 -790 25870 -743
rect 14622 -1071 14668 -790
rect 14880 -831 14926 -790
rect 14880 -1031 15154 -831
rect 14880 -1071 14926 -1031
rect 14622 -1118 14926 -1071
rect 16580 -1118 16976 -790
rect 18356 -1031 18366 -830
rect 18418 -1031 18428 -830
rect 18578 -1031 18588 -831
rect 18640 -1031 18650 -831
rect 20120 -1118 20516 -790
rect 14622 -1276 14668 -1118
rect 14880 -1276 14926 -1118
rect 21870 -1276 21954 -830
rect 22064 -1031 22074 -831
rect 22126 -1031 22136 -831
rect 23641 -1118 24037 -790
rect 25566 -831 25612 -790
rect 25338 -1031 25612 -831
rect 25566 -1071 25612 -1031
rect 25824 -1071 25870 -790
rect 25566 -1118 25870 -1071
rect 25566 -1276 25612 -1118
rect 25824 -1276 25870 -1118
rect 14622 -1323 25870 -1276
rect 14622 -1603 14668 -1323
rect 14880 -1603 14926 -1323
rect 15108 -1602 15154 -1323
rect 15088 -1603 15154 -1602
rect 25566 -1603 25612 -1323
rect 25824 -1603 25870 -1323
rect 14622 -1649 25870 -1603
rect 14622 -1650 15088 -1649
rect 15134 -1650 25870 -1649
rect 21156 -2454 25838 -2408
rect 21156 -2718 21202 -2454
rect 21414 -2718 21460 -2454
rect 25534 -2718 25580 -2454
rect 25792 -2718 25838 -2454
rect 21156 -2764 25838 -2718
rect 21156 -2994 21202 -2764
rect 21414 -2994 21460 -2764
rect 21156 -3040 21231 -2994
rect 21398 -3040 21460 -2994
rect 21156 -3364 21202 -3040
rect 21414 -3364 21460 -3040
rect 21666 -3332 21676 -3072
rect 21728 -3332 21738 -3072
rect 21156 -3410 21218 -3364
rect 21389 -3410 21460 -3364
rect 22341 -3410 22737 -2993
rect 23330 -3332 23340 -3072
rect 23392 -3332 23402 -3072
rect 23592 -3332 23602 -3072
rect 23654 -3332 23664 -3072
rect 21156 -3640 21202 -3410
rect 21414 -3640 21460 -3410
rect 22999 -3481 23186 -3410
rect 23726 -3413 23736 -3361
rect 24073 -3413 24083 -3361
rect 24373 -3410 24769 -2993
rect 25534 -2994 25580 -2764
rect 25792 -2994 25838 -2764
rect 25534 -3040 25604 -2994
rect 25768 -3040 25838 -2994
rect 25256 -3332 25266 -3072
rect 25318 -3332 25328 -3072
rect 25534 -3364 25580 -3040
rect 25792 -3364 25838 -3040
rect 25534 -3410 25600 -3364
rect 25769 -3410 25838 -3364
rect 22999 -3566 23993 -3481
rect 21156 -3686 21221 -3640
rect 21390 -3686 21460 -3640
rect 21156 -4010 21202 -3686
rect 21414 -4010 21460 -3686
rect 21666 -3978 21676 -3718
rect 21728 -3978 21738 -3718
rect 21156 -4056 21230 -4010
rect 21385 -4056 21460 -4010
rect 22336 -4056 22732 -3639
rect 22911 -3689 22921 -3637
rect 23258 -3689 23268 -3637
rect 23806 -3640 23993 -3566
rect 23330 -3978 23340 -3718
rect 23392 -3978 23402 -3718
rect 23592 -3978 23602 -3718
rect 23654 -3978 23664 -3718
rect 24373 -4056 24769 -3639
rect 25534 -3640 25580 -3410
rect 25792 -3640 25838 -3410
rect 25534 -3686 25598 -3640
rect 25766 -3686 25838 -3640
rect 25256 -3978 25266 -3718
rect 25318 -3978 25328 -3718
rect 25534 -4010 25580 -3686
rect 25792 -4010 25838 -3686
rect 25534 -4056 25606 -4010
rect 25764 -4056 25838 -4010
rect 21156 -4286 21202 -4056
rect 21414 -4286 21460 -4056
rect 25534 -4286 25580 -4056
rect 25792 -4286 25838 -4056
rect 21156 -4332 25838 -4286
rect 21156 -4596 21202 -4332
rect 21414 -4596 21460 -4332
rect 25534 -4596 25580 -4332
rect 25792 -4596 25838 -4332
rect 21156 -4642 25838 -4596
<< via1 >>
rect 21788 1989 21840 2189
rect 25338 1989 25390 2189
rect 21788 1458 21840 1657
rect 25338 1456 25390 1657
rect 18366 -499 18418 -299
rect 21852 -499 21904 -299
rect 22074 -499 22126 -299
rect 18366 -1031 18418 -830
rect 18588 -1031 18640 -831
rect 22074 -1031 22126 -831
rect 21676 -3332 21728 -3072
rect 23340 -3332 23392 -3072
rect 23602 -3332 23654 -3072
rect 23736 -3413 24073 -3361
rect 25266 -3332 25318 -3072
rect 21676 -3978 21728 -3718
rect 22921 -3689 23258 -3637
rect 23340 -3978 23392 -3718
rect 23602 -3978 23654 -3718
rect 25266 -3978 25318 -3718
<< metal2 >>
rect 21729 2388 25441 2398
rect 21896 2325 25274 2388
rect 21729 2315 25441 2325
rect 21786 2189 21842 2199
rect 21786 1979 21842 1989
rect 25338 2189 25390 2199
rect 25390 2042 26105 2052
rect 25390 1989 25525 2042
rect 25338 1979 25525 1989
rect 25692 1979 26105 2042
rect 25338 1969 26105 1979
rect 25585 1968 25645 1969
rect 21786 1657 21842 1667
rect 21786 1448 21842 1458
rect 25336 1657 25392 1667
rect 25336 1446 25392 1456
rect 21732 1327 21899 1337
rect 25515 1327 25682 1337
rect 21899 1263 25515 1327
rect 21732 1253 21899 1263
rect 25515 1253 25682 1263
rect 18309 575 22183 585
rect 18476 511 22016 575
rect 18309 501 22183 511
rect 18537 -104 26088 -94
rect 18704 -168 21791 -104
rect 21958 -168 26088 -104
rect 18537 -178 26088 -168
rect 25898 -179 26088 -178
rect 18364 -299 18420 -289
rect 18364 -509 18420 -499
rect 21850 -299 21906 -289
rect 21850 -509 21906 -499
rect 22072 -299 22128 -289
rect 22072 -509 22128 -499
rect 18364 -830 18420 -820
rect 18364 -1041 18420 -1031
rect 18586 -831 18642 -821
rect 18586 -1041 18642 -1031
rect 22072 -831 22128 -821
rect 22072 -1042 22128 -1032
rect 21620 -2847 26121 -2837
rect 21787 -2911 26121 -2847
rect 21620 -2921 26121 -2911
rect 21674 -3072 21730 -3062
rect 21674 -3342 21730 -3332
rect 23338 -3072 23394 -3062
rect 23338 -3342 23394 -3332
rect 23600 -3072 23656 -3062
rect 23600 -3342 23656 -3332
rect 25264 -3072 25320 -3062
rect 25264 -3343 25320 -3333
rect 23736 -3359 24073 -3349
rect 23736 -3425 24073 -3415
rect 23009 -3483 23886 -3482
rect 23009 -3492 23983 -3483
rect 23176 -3493 23983 -3492
rect 23176 -3556 23816 -3493
rect 23009 -3557 23816 -3556
rect 23009 -3566 23983 -3557
rect 23816 -3567 23983 -3566
rect 22921 -3635 23258 -3625
rect 22921 -3701 23258 -3691
rect 21674 -3718 21730 -3708
rect 21674 -3988 21730 -3978
rect 23338 -3718 23394 -3708
rect 23338 -3988 23394 -3978
rect 23600 -3718 23656 -3708
rect 23600 -3988 23656 -3978
rect 25266 -3718 25318 -3708
rect 25318 -3889 26039 -3805
rect 25266 -3988 25318 -3978
rect 21645 -4139 25370 -4129
rect 21645 -4203 21651 -4139
rect 21818 -4203 25203 -4139
rect 21645 -4213 25370 -4203
<< via2 >>
rect 21729 2325 21896 2388
rect 25274 2325 25441 2388
rect 21786 1989 21788 2189
rect 21788 1989 21840 2189
rect 21840 1989 21842 2189
rect 25525 1979 25692 2042
rect 21786 1458 21788 1657
rect 21788 1458 21840 1657
rect 21840 1458 21842 1657
rect 25336 1456 25338 1657
rect 25338 1456 25390 1657
rect 25390 1456 25392 1657
rect 21732 1263 21899 1327
rect 25515 1263 25682 1327
rect 18309 511 18476 575
rect 22016 511 22183 575
rect 18537 -168 18704 -104
rect 21791 -168 21958 -104
rect 18364 -499 18366 -299
rect 18366 -499 18418 -299
rect 18418 -499 18420 -299
rect 21850 -499 21852 -299
rect 21852 -499 21904 -299
rect 21904 -499 21906 -299
rect 22072 -499 22074 -299
rect 22074 -499 22126 -299
rect 22126 -499 22128 -299
rect 18364 -1031 18366 -830
rect 18366 -1031 18418 -830
rect 18418 -1031 18420 -830
rect 18586 -1031 18588 -831
rect 18588 -1031 18640 -831
rect 18640 -1031 18642 -831
rect 22072 -1031 22074 -831
rect 22074 -1031 22126 -831
rect 22126 -1031 22128 -831
rect 22072 -1032 22128 -1031
rect 21620 -2911 21787 -2847
rect 21674 -3332 21676 -3072
rect 21676 -3332 21728 -3072
rect 21728 -3332 21730 -3072
rect 23338 -3332 23340 -3072
rect 23340 -3332 23392 -3072
rect 23392 -3332 23394 -3072
rect 23600 -3332 23602 -3072
rect 23602 -3332 23654 -3072
rect 23654 -3332 23656 -3072
rect 25264 -3332 25266 -3072
rect 25266 -3332 25318 -3072
rect 25318 -3332 25320 -3072
rect 25264 -3333 25320 -3332
rect 23736 -3361 24073 -3359
rect 23736 -3413 24073 -3361
rect 23736 -3415 24073 -3413
rect 23009 -3556 23176 -3492
rect 23816 -3557 23983 -3493
rect 22921 -3637 23258 -3635
rect 22921 -3689 23258 -3637
rect 22921 -3691 23258 -3689
rect 21674 -3978 21676 -3718
rect 21676 -3978 21728 -3718
rect 21728 -3978 21730 -3718
rect 23338 -3978 23340 -3718
rect 23340 -3978 23392 -3718
rect 23392 -3978 23394 -3718
rect 23600 -3978 23602 -3718
rect 23602 -3978 23654 -3718
rect 23654 -3978 23656 -3718
rect 21651 -4203 21818 -4139
rect 25203 -4203 25370 -4139
<< metal3 >>
rect 21719 2388 21906 2393
rect 21719 2325 21729 2388
rect 21896 2325 21906 2388
rect 21719 2320 21906 2325
rect 25264 2388 25451 2393
rect 25264 2325 25274 2388
rect 25441 2325 25451 2388
rect 25264 2320 25451 2325
rect 21776 2189 21852 2320
rect 21776 1989 21786 2189
rect 21842 1989 21852 2189
rect 21776 1984 21852 1989
rect 21776 1657 21852 1662
rect 21776 1458 21786 1657
rect 21842 1458 21852 1657
rect 21776 1332 21852 1458
rect 25326 1657 25402 2320
rect 25515 2042 25702 2047
rect 25515 1979 25525 2042
rect 25692 1979 25702 2042
rect 25515 1974 25702 1979
rect 25326 1456 25336 1657
rect 25392 1456 25402 1657
rect 25326 1451 25402 1456
rect 25583 1332 25647 1974
rect 21722 1327 21909 1332
rect 21722 1263 21732 1327
rect 21899 1263 21909 1327
rect 21722 1258 21909 1263
rect 25505 1327 25692 1332
rect 25505 1263 25515 1327
rect 25682 1263 25692 1327
rect 25505 1258 25692 1263
rect 18299 575 18486 580
rect 18299 511 18309 575
rect 18476 511 18486 575
rect 18299 506 18486 511
rect 22006 575 22193 580
rect 22006 511 22016 575
rect 22183 511 22193 575
rect 22006 506 22193 511
rect 18354 -299 18430 506
rect 18527 -104 18714 -99
rect 18527 -168 18537 -104
rect 18704 -168 18714 -104
rect 18527 -173 18714 -168
rect 21781 -104 21968 -99
rect 21781 -168 21791 -104
rect 21958 -168 21968 -104
rect 21781 -173 21968 -168
rect 18354 -499 18364 -299
rect 18420 -499 18430 -299
rect 18354 -830 18430 -499
rect 18354 -1031 18364 -830
rect 18420 -1031 18430 -830
rect 18354 -1036 18430 -1031
rect 18576 -831 18652 -173
rect 21840 -299 21916 -173
rect 21840 -499 21850 -299
rect 21906 -499 21916 -299
rect 21840 -504 21916 -499
rect 22062 -299 22138 506
rect 22062 -499 22072 -299
rect 22128 -499 22138 -299
rect 18576 -1031 18586 -831
rect 18642 -1031 18652 -831
rect 18576 -1036 18652 -1031
rect 22062 -831 22138 -499
rect 22062 -1032 22072 -831
rect 22128 -1032 22138 -831
rect 22062 -1037 22138 -1032
rect 21610 -2847 21797 -2842
rect 21610 -2911 21620 -2847
rect 21787 -2911 21797 -2847
rect 21610 -2916 21797 -2911
rect 21664 -3072 21740 -2916
rect 21664 -3332 21674 -3072
rect 21730 -3332 21740 -3072
rect 21664 -3337 21740 -3332
rect 23328 -3072 23666 -3067
rect 23328 -3332 23338 -3072
rect 23394 -3332 23600 -3072
rect 23656 -3332 23666 -3072
rect 22999 -3492 23186 -3487
rect 22999 -3556 23009 -3492
rect 23176 -3556 23186 -3492
rect 22999 -3630 23186 -3556
rect 22911 -3635 23268 -3630
rect 22911 -3691 22921 -3635
rect 23258 -3691 23268 -3635
rect 22911 -3696 23268 -3691
rect 21664 -3718 21740 -3713
rect 21664 -3978 21674 -3718
rect 21730 -3978 21740 -3718
rect 21664 -4134 21740 -3978
rect 23328 -3718 23666 -3332
rect 25254 -3072 25330 -3067
rect 25254 -3333 25264 -3072
rect 25320 -3333 25330 -3072
rect 23726 -3359 24083 -3354
rect 23726 -3415 23736 -3359
rect 24073 -3415 24083 -3359
rect 23726 -3420 24083 -3415
rect 23806 -3493 23993 -3420
rect 23806 -3557 23816 -3493
rect 23983 -3557 23993 -3493
rect 23806 -3562 23993 -3557
rect 23328 -3978 23338 -3718
rect 23394 -3978 23600 -3718
rect 23656 -3978 23666 -3718
rect 23328 -3983 23666 -3978
rect 25254 -4134 25330 -3333
rect 21641 -4139 21828 -4134
rect 21641 -4203 21651 -4139
rect 21818 -4203 21828 -4139
rect 21641 -4208 21828 -4203
rect 25193 -4139 25380 -4134
rect 25193 -4203 25203 -4139
rect 25370 -4203 25380 -4139
rect 25193 -4208 25380 -4203
use trans_gate  x1
timestamp 1711994542
transform 1 0 11684 0 1 -1512
box 0 -2380 2272 590
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[0]
timestamp 1712074089
transform 1 0 21460 0 1 2621
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[1]
timestamp 1712074089
transform 1 0 21460 0 1 2089
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[2]
timestamp 1712074089
transform 1 0 21460 0 1 1557
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[3]
timestamp 1712074089
transform 1 0 21460 0 1 1025
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[0]
timestamp 1712242108
transform 1 0 24460 0 1 -3848
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[1]
timestamp 1712242108
transform 1 0 22534 0 1 -3202
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM2[0]
timestamp 1712242108
transform 1 0 24460 0 1 -3202
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM2[1]
timestamp 1712242108
transform 1 0 22534 0 1 -3848
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[0]
timestamp 1712064068
transform -1 0 22646 0 -1 1557
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[1]
timestamp 1712064068
transform 1 0 24532 0 1 2089
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[0]
timestamp 1712150541
transform 1 0 20246 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1712150541
transform 1 0 20246 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[0]
timestamp 1712064068
transform 1 0 24532 0 1 1557
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[1]
timestamp 1712064068
transform 1 0 22646 0 1 2089
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[0]
timestamp 1712150541
transform 1 0 16760 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1712150541
transform 1 0 16760 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[2]
timestamp 1712150541
transform 1 0 23732 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1712150541
transform 1 0 23732 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1711994542
transform 0 1 26587 -1 0 1944
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_L8NDKD  XM8
timestamp 1712242108
transform 0 1 26578 -1 0 -2708
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1711994542
transform 1 0 26564 0 1 175
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1711994542
transform 1 0 26564 0 1 -1094
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1711994542
transform 1 0 18530 0 1 -2538
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1711994542
transform 1 0 18530 0 1 -3052
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1711994542
transform -1 0 20228 0 -1 -3997
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1711994542
transform -1 0 20228 0 -1 -4511
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1711994542
transform 1 0 20414 0 1 1025
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1711994542
transform 1 0 20414 0 1 1557
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1711994542
transform 0 1 26578 -1 0 -4326
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1711994542
transform 1 0 14974 0 1 -2547
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1711994542
transform 1 0 14988 0 1 -3282
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712074089
transform 1 0 25718 0 1 2621
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712074089
transform 1 0 25718 0 1 2089
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712074089
transform 1 0 25718 0 1 1557
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712074089
transform 1 0 25718 0 1 1025
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712074089
transform 1 0 14774 0 1 133
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712074089
transform 1 0 14774 0 1 -399
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712074089
transform 1 0 14774 0 1 -931
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712074089
transform 1 0 14774 0 1 -1463
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712074089
transform 1 0 25718 0 1 133
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712074089
transform 1 0 25718 0 1 -399
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712074089
transform 1 0 25718 0 1 -931
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712074089
transform 1 0 25718 0 1 -1463
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712150541
transform 1 0 16760 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712150541
transform 1 0 20246 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712150541
transform 1 0 23732 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712150541
transform 1 0 16760 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712150541
transform 1 0 20246 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712150541
transform 1 0 23732 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[0]
timestamp 1712064068
transform 1 0 22646 0 1 2621
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[1]
timestamp 1712064068
transform 1 0 24532 0 1 2621
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[2]
timestamp 1712064068
transform 1 0 22646 0 1 1025
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[3]
timestamp 1712064068
transform 1 0 24532 0 1 1025
box -996 -319 996 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712242108
transform 1 0 21308 0 1 -2586
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712242108
transform 1 0 21308 0 1 -4464
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712242108
transform 1 0 25686 0 1 -2586
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712242108
transform 1 0 25686 0 1 -4464
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712242108
transform 1 0 22534 0 1 -2586
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712242108
transform 1 0 24460 0 1 -2586
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[2]
timestamp 1712242108
transform 1 0 22534 0 1 -4464
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[3]
timestamp 1712242108
transform 1 0 24460 0 1 -4464
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712242108
transform 1 0 21308 0 1 -3202
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712242108
transform 1 0 21308 0 1 -3848
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712242108
transform 1 0 25686 0 1 -3202
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712242108
transform 1 0 25686 0 1 -3848
box -328 -388 328 388
<< end >>

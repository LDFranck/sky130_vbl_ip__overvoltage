magic
tech sky130A
timestamp 1713017665
<< pwell >>
rect -164 -179 164 179
<< mvnmos >>
rect -50 -50 50 50
<< mvndiff >>
rect -79 44 -50 50
rect -79 -44 -73 44
rect -56 -44 -50 44
rect -79 -50 -50 -44
rect 50 44 79 50
rect 50 -44 56 44
rect 73 -44 79 44
rect 50 -50 79 -44
<< mvndiffc >>
rect -73 -44 -56 44
rect 56 -44 73 44
<< mvpsubdiff >>
rect -146 155 146 161
rect -146 138 -92 155
rect 92 138 146 155
rect -146 132 146 138
rect -146 107 -117 132
rect -146 -107 -140 107
rect -123 -107 -117 107
rect 117 107 146 132
rect -146 -132 -117 -107
rect 117 -107 123 107
rect 140 -107 146 107
rect 117 -132 146 -107
rect -146 -138 146 -132
rect -146 -155 -92 -138
rect 92 -155 146 -138
rect -146 -161 146 -155
<< mvpsubdiffcont >>
rect -92 138 92 155
rect -140 -107 -123 107
rect 123 -107 140 107
rect -92 -155 92 -138
<< poly >>
rect -50 86 50 94
rect -50 69 -42 86
rect 42 69 50 86
rect -50 50 50 69
rect -50 -69 50 -50
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -50 -94 50 -86
<< polycont >>
rect -42 69 42 86
rect -42 -86 42 -69
<< locali >>
rect -140 138 -92 155
rect 92 138 140 155
rect -140 107 -123 138
rect 123 107 140 138
rect -50 69 -42 86
rect 42 69 50 86
rect -73 44 -56 52
rect -73 -52 -56 -44
rect 56 44 73 52
rect 56 -52 73 -44
rect -50 -86 -42 -69
rect 42 -86 50 -69
rect -140 -138 -123 -107
rect 123 -138 140 -107
rect -140 -155 -92 -138
rect 92 -155 140 -138
<< viali >>
rect -42 69 42 86
rect -73 -44 -56 44
rect 56 -44 73 44
rect -42 -86 42 -69
<< metal1 >>
rect -48 86 48 89
rect -48 69 -42 86
rect 42 69 48 86
rect -48 66 48 69
rect -76 44 -53 50
rect -76 -44 -73 44
rect -56 -44 -53 44
rect -76 -50 -53 -44
rect 53 44 76 50
rect 53 -44 56 44
rect 73 -44 76 44
rect 53 -50 76 -44
rect -48 -69 48 -66
rect -48 -86 -42 -69
rect 42 -86 48 -69
rect -48 -89 48 -86
<< properties >>
string FIXED_BBOX -131 -146 131 146
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1711994542
<< nwell >>
rect 924 144 928 182
rect 1928 144 1932 182
rect 834 90 926 120
rect 918 -1304 920 -1150
<< pwell >>
rect 882 -1870 916 -1716
rect 876 -1874 924 -1870
rect 882 -1880 916 -1874
rect 860 -1892 920 -1880
rect 834 -1922 920 -1892
rect 2108 -2086 2268 -1492
<< mvndiffc >>
rect 882 -1892 916 -1716
<< locali >>
rect 530 500 2272 578
rect 530 380 660 500
rect 2224 380 2272 500
rect 530 286 2272 380
rect 530 144 782 286
rect 924 144 1932 182
rect 2074 144 2268 286
rect 530 -1320 748 144
rect 2108 -1316 2268 144
rect 530 -2080 756 -1494
rect 2108 -2080 2268 -1492
rect 530 -2198 2268 -2080
rect 530 -2318 658 -2198
rect 2222 -2318 2268 -2198
rect 530 -2372 2268 -2318
<< viali >>
rect 660 380 2224 500
rect 882 -1892 916 -1716
rect 658 -2318 2222 -2198
<< metal1 >>
rect 530 500 2272 578
rect 530 380 660 500
rect 2224 380 2272 500
rect 530 286 2272 380
rect 0 0 200 200
rect 1270 140 1280 200
rect 1580 140 1590 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 850 -1088 860 90
rect 916 -1088 926 90
rect 1930 -1088 1940 90
rect 1996 -1088 2006 90
rect 1270 -1200 1280 -1140
rect 1580 -1200 1590 -1140
rect 0 -1600 200 -1400
rect 1270 -1680 1280 -1620
rect 1580 -1680 1590 -1620
rect 0 -2000 200 -1800
rect 850 -1892 860 -1716
rect 916 -1892 926 -1716
rect 1930 -1892 1940 -1716
rect 1996 -1892 2006 -1716
rect 1270 -1992 1280 -1932
rect 1580 -1992 1590 -1932
rect 530 -2198 2268 -2080
rect 530 -2318 658 -2198
rect 2222 -2318 2268 -2198
rect 530 -2372 2268 -2318
<< via1 >>
rect 1280 140 1580 200
rect 860 -1088 916 90
rect 1940 -1088 1996 90
rect 1280 -1200 1580 -1140
rect 1280 -1680 1580 -1620
rect 860 -1892 882 -1716
rect 882 -1892 916 -1716
rect 1940 -1892 1996 -1716
rect 1280 -1992 1580 -1932
<< metal2 >>
rect 1280 200 1580 210
rect 1280 130 1580 140
rect 860 90 916 100
rect 860 -1098 916 -1088
rect 1940 90 1996 100
rect 1940 -1098 1996 -1088
rect 1280 -1140 1580 -1130
rect 1280 -1210 1580 -1200
rect 1280 -1620 1580 -1610
rect 1280 -1690 1580 -1680
rect 860 -1716 916 -1706
rect 860 -1902 916 -1892
rect 1940 -1716 1996 -1706
rect 1940 -1902 1996 -1892
rect 1280 -1932 1580 -1922
rect 1280 -2002 1580 -1992
<< via2 >>
rect 1280 140 1580 200
rect 860 -1088 916 90
rect 1940 -1088 1996 90
rect 1280 -1200 1580 -1140
rect 1280 -1680 1580 -1620
rect 860 -1892 916 -1716
rect 1940 -1892 1996 -1716
rect 1280 -1992 1580 -1932
<< metal3 >>
rect 1280 205 1580 590
rect 1270 200 1590 205
rect 1270 140 1280 200
rect 1580 140 1590 200
rect 1270 135 1590 140
rect 834 90 926 120
rect 834 -1088 860 90
rect 916 -1088 926 90
rect 834 -1093 926 -1088
rect 834 -1304 920 -1093
rect 1280 -1135 1580 135
rect 1926 90 2020 118
rect 1926 -1088 1940 90
rect 1996 -1088 2020 90
rect 1270 -1140 1590 -1135
rect 1270 -1200 1280 -1140
rect 1580 -1200 1590 -1140
rect 1270 -1205 1590 -1200
rect 1926 -1284 2020 -1088
rect 774 -1504 974 -1304
rect 1862 -1484 2062 -1284
rect 834 -1711 920 -1504
rect 1270 -1620 1590 -1615
rect 1270 -1680 1280 -1620
rect 1580 -1680 1590 -1620
rect 1270 -1685 1590 -1680
rect 834 -1716 926 -1711
rect 834 -1892 860 -1716
rect 916 -1892 926 -1716
rect 834 -1897 926 -1892
rect 834 -1922 920 -1897
rect 1280 -1927 1580 -1685
rect 1926 -1716 2020 -1484
rect 1926 -1892 1940 -1716
rect 1996 -1892 2020 -1716
rect 1926 -1926 2020 -1892
rect 1270 -1932 1590 -1927
rect 1270 -1992 1280 -1932
rect 1580 -1992 1590 -1932
rect 1270 -1997 1590 -1992
rect 1280 -2380 1580 -1997
use sky130_fd_pr__nfet_g5v0d10v5_69BJMM  XM1
timestamp 1711651911
transform 1 0 1428 0 1 -1804
box -728 -358 728 358
use sky130_fd_pr__pfet_g5v0d10v5_E7V9VM  XM2
timestamp 1711651911
transform 1 0 1428 0 1 -499
box -758 -897 758 897
<< labels >>
flabel metal1 552 -2372 752 -2172 0 FreeSans 256 0 0 0 vss
port 4 nsew
flabel metal1 532 368 732 568 0 FreeSans 256 0 0 0 avdd
port 3 nsew
flabel metal3 774 -1504 974 -1304 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal3 1862 -1484 2062 -1284 0 FreeSans 256 0 0 0 out
port 5 nsew
flabel metal3 1320 -2380 1520 -2180 0 FreeSans 256 0 0 0 ena
port 2 nsew
flabel metal3 1318 380 1518 580 0 FreeSans 256 0 0 0 ena_b
port 1 nsew
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 in
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 ena_b
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 ena
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 avdd
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 vss
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 out
<< end >>

magic
tech sky130A
timestamp 1712318662
<< pwell >>
rect -514 -179 514 179
<< mvnmos >>
rect -400 -50 400 50
<< mvndiff >>
rect -429 44 -400 50
rect -429 -44 -423 44
rect -406 -44 -400 44
rect -429 -50 -400 -44
rect 400 44 429 50
rect 400 -44 406 44
rect 423 -44 429 44
rect 400 -50 429 -44
<< mvndiffc >>
rect -423 -44 -406 44
rect 406 -44 423 44
<< mvpsubdiff >>
rect -496 155 496 161
rect -496 138 -442 155
rect 442 138 496 155
rect -496 132 496 138
rect -496 107 -467 132
rect -496 -107 -490 107
rect -473 -107 -467 107
rect 467 107 496 132
rect -496 -132 -467 -107
rect 467 -107 473 107
rect 490 -107 496 107
rect 467 -132 496 -107
rect -496 -138 496 -132
rect -496 -155 -442 -138
rect 442 -155 496 -138
rect -496 -161 496 -155
<< mvpsubdiffcont >>
rect -442 138 442 155
rect -490 -107 -473 107
rect 473 -107 490 107
rect -442 -155 442 -138
<< poly >>
rect -400 86 400 94
rect -400 69 -392 86
rect 392 69 400 86
rect -400 50 400 69
rect -400 -69 400 -50
rect -400 -86 -392 -69
rect 392 -86 400 -69
rect -400 -94 400 -86
<< polycont >>
rect -392 69 392 86
rect -392 -86 392 -69
<< locali >>
rect -490 138 -442 155
rect 442 138 490 155
rect -490 107 -473 138
rect 473 107 490 138
rect -400 69 -392 86
rect 392 69 400 86
rect -423 44 -406 52
rect -423 -52 -406 -44
rect 406 44 423 52
rect 406 -52 423 -44
rect -400 -86 -392 -69
rect 392 -86 400 -69
rect -490 -138 -473 -107
rect 473 -138 490 -107
rect -490 -155 -442 -138
rect 442 -155 490 -138
<< viali >>
rect -392 69 392 86
rect -423 -44 -406 44
rect 406 -44 423 44
rect -392 -86 392 -69
<< metal1 >>
rect -398 86 398 89
rect -398 69 -392 86
rect 392 69 398 86
rect -398 66 398 69
rect -426 44 -403 50
rect -426 -44 -423 44
rect -406 -44 -403 44
rect -426 -50 -403 -44
rect 403 44 426 50
rect 403 -44 406 44
rect 423 -44 426 44
rect 403 -50 426 -44
rect -398 -69 398 -66
rect -398 -86 -392 -69
rect 392 -86 398 -69
rect -398 -89 398 -86
<< properties >>
string FIXED_BBOX -481 -146 481 146
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 1 l 8 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

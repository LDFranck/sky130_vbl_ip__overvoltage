magic
tech sky130A
magscale 1 2
timestamp 1712928439
<< pwell >>
rect -183 -7138 183 7138
<< psubdiff >>
rect -147 7068 -51 7102
rect 51 7068 147 7102
rect -147 7006 -113 7068
rect 113 7006 147 7068
rect -147 -7068 -113 -7006
rect 113 -7068 147 -7006
rect -147 -7102 -51 -7068
rect 51 -7102 147 -7068
<< psubdiffcont >>
rect -51 7068 51 7102
rect -147 -7006 -113 7006
rect 113 -7006 147 7006
rect -51 -7102 51 -7068
<< ndiode >>
rect -45 6988 45 7000
rect -45 -6988 -33 6988
rect 33 -6988 45 6988
rect -45 -7000 45 -6988
<< ndiodec >>
rect -33 -6988 33 6988
<< locali >>
rect -147 7068 -51 7102
rect 51 7068 147 7102
rect -147 7006 -113 7068
rect 113 7006 147 7068
rect -33 6988 33 7004
rect -33 -7004 33 -6988
rect -147 -7068 -113 -7006
rect 113 -7068 147 -7006
rect -147 -7102 -51 -7068
rect 51 -7102 147 -7068
<< viali >>
rect -33 -6988 33 6988
<< metal1 >>
rect -39 6988 39 7000
rect -39 -6988 -33 6988
rect 33 -6988 39 6988
rect -39 -7000 39 -6988
<< properties >>
string FIXED_BBOX -130 -7085 130 7085
string gencell sky130_fd_pr__diode_pw2nd_05v5
string library sky130
string parameters w 0.45 l 70 area 31.5 peri 140.9 nx 1 ny 1 dummy 0 lmin 0.45 wmin 0.45 elc 1 erc 1 etc 1 ebc 1 doverlap 0 compatible {sky130_fd_pr__diode_pw2nd_05v5 sky130_fd_pr__diode_pw2nd_05v5_lvt  sky130_fd_pr__diode_pw2nd_05v5_nvt sky130_fd_pr__diode_pw2nd_11v0} full_metal 1 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

* expanding   symbol:  sky130_vbl_ip__overvoltage.sym # of pins=11
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/sky130_vbl_ip__overvoltage.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/sky130_vbl_ip__overvoltage.sch
.subckt sky130_vbl_ip__overvoltage avdd dvdd ena vtrip[3] vss ibias vtrip[2] ovout vbg vtrip[1] vtrip[0]
*.iopin avdd
*.iopin dvdd
*.ipin ena
*.iopin vss
*.ipin vtrip[3]
*.opin ovout
*.ipin vbg
*.ipin vtrip[2]
*.ipin vtrip[1]
*.ipin vtrip[0]
*.ipin ibias
x1 avdd dvdd net1 vtrip[3] A NotA vss LevelShifter
XVBIAS1 avdd net1 ena vss halfvdd_vbias
x2 avdd dvdd net1 vtrip[2] B NotB vss LevelShifter
x3 avdd dvdd net1 vtrip[1] C NotC vss LevelShifter
x4 avdd dvdd net1 vtrip[0] D NotD vss LevelShifter
x5 net4 net5 net6 net7 net8 net9 net10 avdd vss net11 A NotA B NotB C net2 NotC D NotD net3 net12 net13 net14 net15 net16 net17
+ net18 DemuxCompleto
x6 avdd net4 net5 net6 net7 net8 net9 net10 net11 net3 net12 net13 net14 net15 net16 net17 net18 vss ena divisor_completo
x7 dvdd ovout vbg net2 ena ibias vss comp_hyst
.ends


* expanding   symbol:  LevelShifter.sym # of pins=7
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/LevelShifter.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/LevelShifter.sch
.subckt LevelShifter avdd dvdd bias in out out_b vss
*.ipin in
*.iopin dvdd
*.opin out
*.opin out_b
*.iopin avdd
*.ipin bias
*.iopin vss
XM3 out in_b vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 in_b in dvdd dvdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net1 net2 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net2 net1 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 out_b bias net1 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 out bias net2 avdd sky130_fd_pr__pfet_g5v0d10v5 L=1 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 out_b in vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 in_b in vss vss sky130_fd_pr__nfet_g5v0d10v5 L=1 W=10 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  halfvdd_vbias.sym # of pins=4
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/halfvdd_vbias.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/halfvdd_vbias.sch
.subckt halfvdd_vbias avdd bias ena vss
*.ipin ena
*.iopin vss
*.iopin avdd
*.opin bias
XM1 net3 net3 avdd avdd sky130_fd_pr__pfet_g5v0d10v5 L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 net3 bias bias sky130_fd_pr__pfet_g5v0d10v5 L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net2 bias bias sky130_fd_pr__pfet_g5v0d10v5 L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net2 net1 net1 sky130_fd_pr__pfet_g5v0d10v5 L=10 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 ena vss vss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  DemuxCompleto.sym # of pins=27
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/DemuxCompleto.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/DemuxCompleto.sch
.subckt DemuxCompleto in_0000 in_0001 in_0010 in_0011 in_0100 in_0101 in_0110 avdd vss in_0111 vtrip_3 vtrip_3_b vtrip_2 vtrip_2_b
+ vtrip_1 out vtrip_1_b vtrip_0 vtrip_0_b in_1000 in_1001 in_1010 in_1011 in_1100 in_1101 in_1110 in_1111
*.ipin in_0000
*.ipin in_0001
*.ipin in_0010
*.ipin in_0011
*.ipin in_0100
*.ipin in_0101
*.ipin in_0110
*.ipin in_0111
*.ipin in_1000
*.ipin in_1001
*.ipin in_1010
*.ipin in_1011
*.ipin in_1110
*.ipin in_1111
*.ipin in_1100
*.ipin in_1101
*.opin out
*.ipin vtrip_3
*.ipin vtrip_3_b
*.ipin vtrip_2
*.ipin vtrip_2_b
*.ipin vtrip_1
*.ipin vtrip_1_b
*.ipin vtrip_0
*.ipin vtrip_0_b
*.iopin avdd
*.iopin vss
x1 vtrip_3 avdd net5 out vss vtrip_3_b T_gate
x2 vtrip_3_b avdd net6 out vss vtrip_3 T_gate
x3 vtrip_2 avdd net2 net6 vss vtrip_2_b T_gate
x4 vtrip_2_b avdd net4 net5 vss vtrip_2 T_gate
x5 vtrip_2_b avdd net3 net6 vss vtrip_2 T_gate
x6 vtrip_2 avdd net1 net5 vss vtrip_2_b T_gate
x7 vtrip_1 avdd net7 net1 vss vtrip_1_b T_gate
x8 vtrip_1_b avdd net8 net1 vss vtrip_1 T_gate
x9 vtrip_1 avdd net9 net4 vss vtrip_1_b T_gate
x10 vtrip_1_b avdd net10 net4 vss vtrip_1 T_gate
x11 vtrip_1 avdd net11 net2 vss vtrip_1_b T_gate
x12 vtrip_1_b avdd net12 net2 vss vtrip_1 T_gate
x13 vtrip_1 avdd net13 net3 vss vtrip_1_b T_gate
x14 vtrip_1_b avdd net14 net3 vss vtrip_1 T_gate
x15 vtrip_0 avdd in_0000 net7 vss vtrip_0_b T_gate
x16 vtrip_0_b avdd in_0001 net7 vss vtrip_0 T_gate
x17 vtrip_0 avdd in_0010 net8 vss vtrip_0_b T_gate
x18 vtrip_0_b avdd in_0011 net8 vss vtrip_0 T_gate
x19 vtrip_0 avdd in_0100 net9 vss vtrip_0_b T_gate
x20 vtrip_0_b avdd in_0101 net9 vss vtrip_0 T_gate
x21 vtrip_0 avdd in_0110 net10 vss vtrip_0_b T_gate
x22 vtrip_0_b avdd in_0111 net10 vss vtrip_0 T_gate
x23 vtrip_0 avdd in_1000 net11 vss vtrip_0_b T_gate
x24 vtrip_0_b avdd in_1001 net11 vss vtrip_0 T_gate
x25 vtrip_0 avdd in_1010 net12 vss vtrip_0_b T_gate
x26 vtrip_0_b avdd in_1011 net12 vss vtrip_0 T_gate
x27 vtrip_0 avdd in_1100 net13 vss vtrip_0_b T_gate
x28 vtrip_0_b avdd in_1101 net15 vss vtrip_0 T_gate
x29 vtrip_0 avdd in_1110 net14 vss vtrip_0_b T_gate
x30 vtrip_0_b avdd in_1111 net14 vss vtrip_0 T_gate
.ends


* expanding   symbol:  divisor_completo.sym # of pins=19
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/divisor_completo.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/divisor_completo.sch
.subckt divisor_completo avdd out_0000 out_0001 out_0010 out_0011 out_0100 out_0101 out_0110 out_0111 out_1000 out_1001 out_1010
+ out_1011 out_1100 out_1101 out_1110 out_1111 vss ena
*.ipin ena
*.iopin vss
*.iopin avdd
*.opin out_1110
*.opin out_1101
*.opin out_1100
*.opin out_1011
*.opin out_1010
*.opin out_1001
*.opin out_1000
*.opin out_0000
*.opin out_0001
*.opin out_0010
*.opin out_0011
*.opin out_0100
*.opin out_0101
*.opin out_0110
*.opin out_0111
*.opin out_1111
x1 out_0000 out_0001 vss div_voltage
x2 out_0001 out_0010 vss div_voltage
x3 out_0010 out_0011 vss div_voltage
x4 out_0011 out_0100 vss div_voltage
x5 out_0100 out_0101 vss div_voltage
x6 out_0101 out_0110 vss div_voltage
x7 out_0110 out_0111 vss div_voltage
x8 out_0111 out_1000 vss div_voltage
x9 out_1000 out_1001 vss div_voltage
x10 out_1001 out_1010 vss div_voltage
x11 out_1010 out_1011 vss div_voltage
x12 out_1011 out_1100 vss div_voltage
x13 out_1100 out_1101 vss div_voltage
x14 out_1101 out_1110 vss div_voltage
x15 out_1110 out_1111 vss div_voltage
XR1 out_0000 avdd vss sky130_fd_pr__res_xhigh_po_0p35 L=92.4 mult=1 m=1
XR2 net1 out_1111 vss sky130_fd_pr__res_xhigh_po_0p35 L=30.1 mult=1 m=1
XM1 net1 ena vss vss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=5 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  comp_hyst.sym # of pins=7
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/comp_hyst.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/comp_hyst.sch
.subckt comp_hyst dvdd out - + ena ibias vss
*.iopin dvdd
*.ipin -
*.ipin +
*.opin out
*.ipin ibias
*.ipin ena
*.iopin vss
XM4 net3 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 ena dvdd dvdd sky130_fd_pr__pfet_01v8 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net3 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net1 net3 dvdd dvdd sky130_fd_pr__pfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM10 net2 net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 ibias ibias vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 vx ibias vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2[0] out net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2[1] out net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2[2] out net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2[3] out net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13[0] out net1 vss vss sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13[1] out net1 vss vss sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13[2] out net1 vss vss sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13[3] out net1 vss vss sky130_fd_pr__nfet_01v8 L=1 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM20 out ena_b vss vss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3[0] net3 - vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3[1] net3 - vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3[2] net3 - vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3[3] net3 - vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4[0] net2 + vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4[1] net2 + vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4[2] net2 + vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4[3] net2 + vx vss sky130_fd_pr__nfet_g5v0d10v5 L=10 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 ibias ena_b vss vss sky130_fd_pr__nfet_01v8 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1[0] net3 net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1[1] net3 net2 dvdd dvdd sky130_fd_pr__pfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 ena_b ena vss vss sky130_fd_pr__nfet_g5v0d10v5 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 ena_b ena dvdd dvdd sky130_fd_pr__pfet_g5v0d10v5 L=3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 net1 vss vss sky130_fd_pr__nfet_01v8 L=20 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  T_gate.sym # of pins=6
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/T_gate.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/T_gate.sch
.subckt T_gate vtrip avdd in out vss vtrip_b
*.iopin avdd
*.iopin vss
*.ipin vtrip
*.ipin vtrip_b
*.ipin in
*.opin out
XM1 in vtrip_b out vss sky130_fd_pr__nfet_g5v0d10v5 L=5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 in vtrip out avdd sky130_fd_pr__pfet_g5v0d10v5 L=5 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  div_voltage.sym # of pins=3
** sym_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/div_voltage.sym
** sch_path: /home/vblabs/Music/sky130_vbl_ip__overvoltage/xschem/div_voltage.sch
.subckt div_voltage v1 v2 vss
*.iopin vss
*.iopin v1
*.iopin v2
XR1 net1 v1 vss sky130_fd_pr__res_xhigh_po_0p35 L=0.70 mult=1 m=1
XR2 v2 net1 vss sky130_fd_pr__res_xhigh_po_0p35 L=0.70 mult=1 m=1
.ends

.GLOBAL GND
.end

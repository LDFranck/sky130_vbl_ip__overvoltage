magic
tech sky130A
magscale 1 2
timestamp 1712171732
<< nwell >>
rect 21566 838 21612 2808
rect 21776 2194 21852 2323
rect 23565 2189 23612 2434
rect 25180 2315 25274 2398
rect 25390 2024 25526 2052
rect 25338 1969 25525 1982
rect 25583 1972 25585 1974
rect 25645 1972 25647 1974
rect 25326 1662 25402 1865
rect 21776 1263 21852 1453
rect 14622 273 14854 320
rect 14622 -7 14668 273
rect 14880 -7 14926 273
rect 15108 -7 15154 287
rect 25807 273 25870 320
rect 14622 -55 14926 -7
rect 15090 -22 15154 -7
rect 15090 -26 15151 -22
rect 15090 -54 15108 -26
rect 14622 -211 14668 -55
rect 14880 -211 14926 -55
rect 14622 -258 14926 -211
rect 14622 -539 14668 -258
rect 14880 -299 14926 -258
rect 25566 -211 25612 273
rect 25824 -7 25870 273
rect 25802 -54 25870 -7
rect 25824 -211 25870 -54
rect 25566 -258 25870 -211
rect 25566 -299 25612 -258
rect 14880 -499 15108 -299
rect 25338 -499 25612 -299
rect 14880 -539 14926 -499
rect 14622 -586 14926 -539
rect 14622 -743 14668 -586
rect 14880 -743 14926 -586
rect 14622 -790 14926 -743
rect 14622 -1071 14668 -790
rect 14880 -831 14926 -790
rect 25566 -539 25612 -499
rect 25824 -539 25870 -258
rect 25566 -586 25870 -539
rect 25566 -743 25612 -586
rect 25824 -743 25870 -586
rect 25566 -790 25870 -743
rect 25566 -831 25612 -790
rect 14880 -1031 15108 -831
rect 25338 -1031 25612 -831
rect 14880 -1071 14926 -1031
rect 14622 -1118 14926 -1071
rect 14622 -1276 14668 -1118
rect 14880 -1276 14926 -1118
rect 25566 -1071 25612 -1031
rect 25824 -1071 25870 -790
rect 25566 -1118 25870 -1071
rect 25566 -1276 25612 -1118
rect 25824 -1276 25870 -1118
rect 14622 -1323 14926 -1276
rect 15085 -1308 15108 -1276
rect 15085 -1321 15152 -1308
rect 15085 -1323 15154 -1321
rect 14622 -1603 14668 -1323
rect 14880 -1603 14926 -1323
rect 14622 -1650 14926 -1603
rect 15108 -1625 15154 -1323
rect 15134 -1626 15154 -1625
rect 25566 -1323 25870 -1276
rect 25566 -1603 25612 -1323
rect 25824 -1603 25870 -1323
rect 25566 -1650 25870 -1603
<< poly >>
rect 25645 1972 25647 1974
<< metal1 >>
rect 21308 2762 25871 2808
rect 21308 2480 21354 2762
rect 21566 2480 21612 2762
rect 21794 2480 21841 2762
rect 23452 2480 23499 2762
rect 23680 2480 23727 2762
rect 25339 2480 25386 2762
rect 25566 2480 25612 2762
rect 25825 2480 25871 2762
rect 21308 2434 25871 2480
rect 21308 2276 21354 2434
rect 21566 2276 21612 2434
rect 21308 2230 21612 2276
rect 21308 1948 21354 2230
rect 21566 1948 21612 2230
rect 21778 1989 21788 2189
rect 21840 1989 21850 2189
rect 22418 1948 22815 2277
rect 23565 2189 23612 2434
rect 23453 1989 23726 2189
rect 24340 1948 24737 2277
rect 25566 2276 25612 2434
rect 25825 2276 25871 2434
rect 25566 2230 25871 2276
rect 25328 1989 25338 2189
rect 25390 1989 25400 2189
rect 25566 1948 25612 2230
rect 25825 1948 25871 2230
rect 21308 1902 21612 1948
rect 21308 1744 21354 1902
rect 21566 1744 21612 1902
rect 21308 1698 21612 1744
rect 21850 1698 25327 1948
rect 25566 1902 25871 1948
rect 25566 1744 25612 1902
rect 25825 1744 25871 1902
rect 25566 1698 25871 1744
rect 21308 1416 21354 1698
rect 21566 1416 21612 1698
rect 21778 1458 21788 1657
rect 21840 1458 21850 1657
rect 21308 1370 21612 1416
rect 21308 1212 21354 1370
rect 21566 1212 21612 1370
rect 22418 1369 22815 1698
rect 23451 1457 23726 1657
rect 23565 1212 23612 1457
rect 24339 1370 24736 1698
rect 25328 1456 25338 1657
rect 25390 1456 25400 1657
rect 25566 1416 25612 1698
rect 25825 1416 25871 1698
rect 25566 1370 25871 1416
rect 25566 1212 25612 1370
rect 25825 1212 25871 1370
rect 21308 1166 25871 1212
rect 21308 884 21354 1166
rect 21566 884 21612 1166
rect 21794 884 21841 1166
rect 23452 884 23499 1166
rect 23680 884 23727 1166
rect 25338 884 25385 1166
rect 25566 884 25612 1166
rect 25825 884 25871 1166
rect 21308 838 25871 884
rect 14622 273 25870 320
rect 14622 -7 14668 273
rect 14880 -7 14926 273
rect 15108 -7 15154 273
rect 25566 -7 25612 273
rect 25824 -7 25870 273
rect 14622 -54 25870 -7
rect 14622 -55 14926 -54
rect 14622 -211 14668 -55
rect 14880 -211 14926 -55
rect 14622 -258 14926 -211
rect 14622 -539 14668 -258
rect 14880 -299 14926 -258
rect 14880 -499 15154 -299
rect 14880 -539 14926 -499
rect 14622 -586 14926 -539
rect 16580 -540 16976 -211
rect 20120 -540 20516 -210
rect 23640 -540 24036 -210
rect 25566 -211 25612 -54
rect 25824 -211 25870 -54
rect 25566 -258 25870 -211
rect 25566 -299 25612 -258
rect 25338 -499 25612 -299
rect 25566 -539 25612 -499
rect 25824 -539 25870 -258
rect 14622 -743 14668 -586
rect 14880 -743 14926 -586
rect 14622 -790 14926 -743
rect 15164 -790 25328 -540
rect 25566 -586 25870 -539
rect 25566 -743 25612 -586
rect 25824 -743 25870 -586
rect 25566 -790 25870 -743
rect 14622 -1071 14668 -790
rect 14880 -831 14926 -790
rect 14880 -1031 15154 -831
rect 14880 -1071 14926 -1031
rect 14622 -1118 14926 -1071
rect 16580 -1118 16976 -790
rect 20120 -1118 20516 -790
rect 23641 -1118 24037 -790
rect 25566 -831 25612 -790
rect 25338 -1031 25612 -831
rect 25566 -1071 25612 -1031
rect 25824 -1071 25870 -790
rect 25566 -1118 25870 -1071
rect 14622 -1276 14668 -1118
rect 14880 -1276 14926 -1118
rect 25566 -1276 25612 -1118
rect 25824 -1276 25870 -1118
rect 14622 -1323 25870 -1276
rect 14622 -1603 14668 -1323
rect 14880 -1603 14926 -1323
rect 15108 -1602 15154 -1323
rect 15088 -1603 15154 -1602
rect 25566 -1603 25612 -1323
rect 25824 -1603 25870 -1323
rect 14622 -1649 25870 -1603
rect 14622 -1650 15088 -1649
rect 15134 -1650 25870 -1649
<< via1 >>
rect 21788 1989 21840 2189
rect 25338 1989 25390 2189
rect 21788 1458 21840 1657
rect 25338 1456 25390 1657
<< metal2 >>
rect 21729 2388 25441 2398
rect 21896 2325 25274 2388
rect 21729 2315 25441 2325
rect 21786 2189 21842 2199
rect 21786 1979 21842 1989
rect 25338 2189 25390 2199
rect 25390 2042 26105 2052
rect 25390 1989 25525 2042
rect 25338 1979 25525 1989
rect 25692 1979 26105 2042
rect 25338 1969 26105 1979
rect 25585 1968 25645 1969
rect 21786 1657 21842 1667
rect 21786 1448 21842 1458
rect 25336 1657 25392 1667
rect 25336 1446 25392 1456
rect 21732 1327 21899 1337
rect 25515 1327 25682 1337
rect 21899 1263 25515 1327
rect 21732 1253 21899 1263
rect 25515 1253 25682 1263
<< via2 >>
rect 21729 2325 21896 2388
rect 25274 2325 25441 2388
rect 21786 1989 21788 2189
rect 21788 1989 21840 2189
rect 21840 1989 21842 2189
rect 25525 1979 25692 2042
rect 21786 1458 21788 1657
rect 21788 1458 21840 1657
rect 21840 1458 21842 1657
rect 25336 1456 25338 1657
rect 25338 1456 25390 1657
rect 25390 1456 25392 1657
rect 21732 1263 21899 1327
rect 25515 1263 25682 1327
<< metal3 >>
rect 21719 2388 21906 2393
rect 21719 2325 21729 2388
rect 21896 2325 21906 2388
rect 21719 2320 21906 2325
rect 25264 2388 25451 2393
rect 25264 2325 25274 2388
rect 25441 2325 25451 2388
rect 25264 2320 25451 2325
rect 21776 2189 21852 2320
rect 21776 1989 21786 2189
rect 21842 1989 21852 2189
rect 21776 1984 21852 1989
rect 21776 1657 21852 1662
rect 21776 1458 21786 1657
rect 21842 1458 21852 1657
rect 21776 1332 21852 1458
rect 25326 1657 25402 2320
rect 25515 2042 25702 2047
rect 25515 1979 25525 2042
rect 25692 1979 25702 2042
rect 25515 1974 25702 1979
rect 25326 1456 25336 1657
rect 25392 1456 25402 1657
rect 25326 1451 25402 1456
rect 25583 1332 25647 1974
rect 21722 1327 21909 1332
rect 21722 1263 21732 1327
rect 21899 1263 21909 1327
rect 21722 1258 21909 1263
rect 25505 1327 25692 1332
rect 25505 1263 25515 1327
rect 25682 1263 25692 1327
rect 25505 1258 25692 1263
use trans_gate  x1
timestamp 1711994542
transform 1 0 10405 0 1 -914
box 0 -2380 2272 590
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[0]
timestamp 1712074089
transform 1 0 21460 0 1 2621
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[1]
timestamp 1712074089
transform 1 0 21460 0 1 2089
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[2]
timestamp 1712074089
transform 1 0 21460 0 1 1557
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[3]
timestamp 1712074089
transform 1 0 21460 0 1 1025
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[0]
timestamp 1712150472
transform 1 0 24460 0 1 -3608
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[1]
timestamp 1712150472
transform 1 0 22534 0 1 -2962
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM2[0]
timestamp 1712150472
transform 1 0 24460 0 1 -2962
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM2[1]
timestamp 1712150472
transform 1 0 22534 0 1 -3608
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[0]
timestamp 1712064068
transform -1 0 22646 0 -1 1557
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[1]
timestamp 1712064068
transform 1 0 24532 0 1 2089
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[0]
timestamp 1712150541
transform 1 0 20246 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1712150541
transform 1 0 20246 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[0]
timestamp 1712064068
transform 1 0 24532 0 1 1557
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[1]
timestamp 1712064068
transform 1 0 22646 0 1 2089
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[0]
timestamp 1712150541
transform 1 0 16760 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1712150541
transform 1 0 16760 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[2]
timestamp 1712150541
transform 1 0 23732 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1712150541
transform 1 0 23732 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1711994542
transform 0 1 26589 -1 0 506
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_697RXD  XM8
timestamp 1711994542
transform 0 1 26570 -1 0 -4082
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1711994542
transform 1 0 26564 0 1 -1263
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1711994542
transform 1 0 26564 0 1 -2498
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1711994542
transform 1 0 18530 0 1 -2298
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1711994542
transform 1 0 18530 0 1 -2812
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1711994542
transform -1 0 20228 0 -1 -3757
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1711994542
transform -1 0 20228 0 -1 -4271
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1711994542
transform 1 0 20414 0 1 1025
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1711994542
transform 1 0 20414 0 1 1557
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1711994542
transform 1 0 25519 0 1 -5021
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1711994542
transform 1 0 13727 0 1 -1463
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1711994542
transform 1 0 13727 0 1 -2298
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712074089
transform 1 0 25718 0 1 2621
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712074089
transform 1 0 25718 0 1 2089
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712074089
transform 1 0 25718 0 1 1557
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712074089
transform 1 0 25718 0 1 1025
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712074089
transform 1 0 14774 0 1 133
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712074089
transform 1 0 14774 0 1 -399
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712074089
transform 1 0 14774 0 1 -931
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712074089
transform 1 0 14774 0 1 -1463
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712074089
transform 1 0 25718 0 1 133
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712074089
transform 1 0 25718 0 1 -399
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712074089
transform 1 0 25718 0 1 -931
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712074089
transform 1 0 25718 0 1 -1463
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712150541
transform 1 0 16760 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712150541
transform 1 0 20246 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712150541
transform 1 0 23732 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712150541
transform 1 0 16760 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712150541
transform 1 0 20246 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712150541
transform 1 0 23732 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[0]
timestamp 1712064068
transform 1 0 22646 0 1 2621
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[1]
timestamp 1712064068
transform 1 0 24532 0 1 2621
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[2]
timestamp 1712064068
transform 1 0 22646 0 1 1025
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[3]
timestamp 1712064068
transform 1 0 24532 0 1 1025
box -996 -319 996 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712151124
transform 1 0 21308 0 1 -2346
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712151124
transform 1 0 21308 0 1 -4224
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712151124
transform 1 0 25686 0 1 -2346
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712151124
transform 1 0 25686 0 1 -4224
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712150472
transform 1 0 22534 0 1 -2346
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712150472
transform 1 0 24460 0 1 -2346
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[2]
timestamp 1712150472
transform 1 0 22534 0 1 -4224
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[3]
timestamp 1712150472
transform 1 0 24460 0 1 -4224
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712151124
transform 1 0 21308 0 1 -2962
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712151124
transform 1 0 21308 0 1 -3608
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712151124
transform 1 0 25686 0 1 -2962
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712151124
transform 1 0 25686 0 1 -3608
box -328 -388 328 388
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712947935
<< locali >>
rect 1298 510 2658 522
rect 1298 442 1315 510
rect 2641 442 2658 510
rect 1298 430 2658 442
rect 1295 -2016 2655 -2004
rect 1295 -2084 1312 -2016
rect 2638 -2084 2655 -2016
rect 1295 -2096 2655 -2084
<< viali >>
rect 1315 442 2641 510
rect 1312 -2084 2638 -2016
<< metal1 >>
rect 1298 510 2658 522
rect 1298 442 1315 510
rect 2641 442 2658 510
rect 1298 430 2658 442
rect 1468 259 1478 311
rect 2478 259 2488 311
rect 1410 -989 1420 211
rect 1472 -989 1482 211
rect 2513 -986 2573 211
rect 1468 -1089 1478 -1037
rect 2478 -1089 2488 -1037
rect 2516 -1273 2573 -986
rect 1296 -1349 2573 -1273
rect 1373 -1594 1437 -1349
rect 1465 -1546 1475 -1494
rect 2475 -1546 2485 -1494
rect 1373 -1794 1469 -1594
rect 2471 -1794 2481 -1594
rect 2533 -1794 2543 -1594
rect 1465 -1894 1475 -1842
rect 2475 -1894 2485 -1842
rect 1295 -2016 2655 -2004
rect 1295 -2084 1312 -2016
rect 2638 -2084 2655 -2016
rect 1295 -2096 2655 -2084
<< via1 >>
rect 1478 259 2478 311
rect 1420 -989 1472 211
rect 1478 -1089 2478 -1037
rect 1475 -1546 2475 -1494
rect 2481 -1794 2533 -1594
rect 1475 -1894 2475 -1842
<< metal2 >>
rect 1478 315 2658 325
rect 1478 311 2508 315
rect 2478 259 2508 311
rect 2648 259 2658 315
rect 1478 249 2658 259
rect 1418 211 1474 221
rect 1418 -999 1474 -989
rect 1478 -1037 2658 -1027
rect 2478 -1089 2508 -1037
rect 1478 -1093 2508 -1089
rect 2648 -1093 2658 -1037
rect 1478 -1103 2658 -1093
rect 1373 -1283 2655 -1273
rect 1513 -1339 2433 -1283
rect 2573 -1339 2655 -1283
rect 1373 -1349 2655 -1339
rect 1247 -1490 2475 -1480
rect 1247 -1546 1259 -1490
rect 1399 -1494 2475 -1490
rect 1399 -1546 1475 -1494
rect 1247 -1556 2475 -1546
rect 2479 -1594 2535 -1584
rect 2479 -1804 2535 -1794
rect 1247 -1842 2475 -1832
rect 1247 -1898 1259 -1842
rect 1399 -1894 1475 -1842
rect 1399 -1898 2475 -1894
rect 1247 -1908 2475 -1898
<< via2 >>
rect 2508 259 2648 315
rect 1418 -989 1420 211
rect 1420 -989 1472 211
rect 1472 -989 1474 211
rect 2508 -1093 2648 -1037
rect 1373 -1339 1513 -1283
rect 2433 -1339 2573 -1283
rect 1259 -1546 1399 -1490
rect 2479 -1794 2481 -1594
rect 2481 -1794 2533 -1594
rect 2533 -1794 2535 -1594
rect 1259 -1898 1399 -1842
<< metal3 >>
rect 2498 315 2658 325
rect 2498 259 2508 315
rect 2648 259 2658 315
rect 1408 211 1484 216
rect 1408 -989 1418 211
rect 1474 -989 1484 211
rect 1408 -1278 1484 -989
rect 2498 -1037 2658 259
rect 2498 -1093 2508 -1037
rect 2648 -1093 2658 -1037
rect 2498 -1098 2658 -1093
rect 1363 -1283 1523 -1278
rect 1363 -1339 1373 -1283
rect 1513 -1339 1523 -1283
rect 1363 -1344 1523 -1339
rect 2423 -1283 2583 -1278
rect 2423 -1339 2433 -1283
rect 2573 -1339 2583 -1283
rect 2423 -1344 2583 -1339
rect 1247 -1490 1409 -1480
rect 1247 -1546 1259 -1490
rect 1399 -1546 1409 -1490
rect 1247 -1842 1409 -1546
rect 2469 -1594 2545 -1344
rect 2469 -1794 2479 -1594
rect 2535 -1794 2545 -1594
rect 2469 -1799 2545 -1794
rect 1247 -1898 1259 -1842
rect 1399 -1898 1409 -1842
rect 1247 -1908 1409 -1898
use sky130_fd_pr__nfet_g5v0d10v5_69BJMM  XM1
timestamp 1712777902
transform 1 0 1975 0 1 -1694
box -728 -358 728 358
use sky130_fd_pr__pfet_g5v0d10v5_E7V9VM  XM2
timestamp 1712777902
transform 1 0 1978 0 1 -389
box -758 -897 758 897
<< labels >>
flabel metal2 2573 -1349 2655 -1273 0 FreeSans 640 0 0 0 out
port 6 nsew
flabel metal1 1296 -1349 1373 -1273 0 FreeSans 640 0 0 0 in
port 1 nsew
flabel metal3 1247 -1908 1409 -1832 0 FreeSans 640 0 0 0 ena
port 3 nsew
flabel metal3 2498 249 2658 325 0 FreeSans 640 0 0 0 ena_b
port 2 nsew
flabel metal1 1295 -2096 2655 -2004 0 FreeSans 1280 0 0 0 vss
port 5 nsew
flabel metal1 1298 430 2658 522 0 FreeSans 1280 0 0 0 avdd
port 4 nsew
<< end >>

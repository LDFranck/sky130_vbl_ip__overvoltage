magic
tech sky130A
magscale 1 2
timestamp 1712319635
<< nwell >>
rect 25583 1972 25585 1974
rect 25645 1972 25647 1974
rect 25326 1662 25402 1865
rect 15090 -22 15108 -7
rect 15090 -26 15151 -22
rect 15090 -54 15108 -26
rect 14668 -1650 14880 -1603
<< poly >>
rect 25645 1972 25647 1974
<< metal1 >>
rect 21308 2762 25871 2808
rect 21308 2480 21354 2762
rect 21566 2480 21612 2762
rect 21794 2480 21841 2762
rect 23452 2480 23499 2762
rect 23680 2480 23727 2762
rect 25339 2480 25386 2762
rect 25566 2480 25612 2762
rect 25825 2480 25871 2762
rect 21308 2434 25871 2480
rect 21308 2276 21354 2434
rect 21566 2276 21612 2434
rect 21308 2230 21612 2276
rect 21308 1948 21354 2230
rect 21566 1948 21612 2230
rect 21778 1989 21788 2189
rect 21840 1989 21850 2189
rect 22418 1948 22815 2277
rect 23504 2189 23673 2434
rect 23453 1989 23726 2189
rect 24340 1948 24737 2277
rect 25566 2276 25612 2434
rect 25825 2276 25871 2434
rect 25566 2230 25871 2276
rect 25328 1989 25338 2189
rect 25390 1989 25400 2189
rect 25566 1948 25612 2230
rect 25825 1948 25871 2230
rect 21308 1902 21612 1948
rect 21308 1744 21354 1902
rect 21566 1744 21612 1902
rect 21308 1698 21612 1744
rect 21850 1698 25327 1948
rect 25566 1902 25871 1948
rect 25566 1744 25612 1902
rect 25825 1744 25871 1902
rect 25566 1698 25871 1744
rect 21308 1416 21354 1698
rect 21566 1416 21612 1698
rect 21778 1458 21788 1657
rect 21840 1458 21850 1657
rect 21308 1370 21612 1416
rect 21308 1212 21354 1370
rect 21566 1212 21612 1370
rect 22418 1369 22815 1698
rect 23451 1457 23726 1657
rect 23499 1212 23668 1457
rect 24339 1370 24736 1698
rect 25328 1456 25338 1657
rect 25390 1456 25400 1657
rect 25566 1416 25612 1698
rect 25825 1416 25871 1698
rect 25566 1370 25871 1416
rect 25566 1212 25612 1370
rect 25825 1212 25871 1370
rect 21308 1166 25871 1212
rect 21308 884 21354 1166
rect 21566 884 21612 1166
rect 21794 884 21841 1166
rect 23452 884 23499 1166
rect 23680 884 23727 1166
rect 25338 884 25385 1166
rect 25566 884 25612 1166
rect 25825 884 25871 1166
rect 21308 838 25871 884
rect 14622 273 25870 320
rect 14622 -7 14668 273
rect 14880 -7 14926 273
rect 15108 -7 15154 273
rect 25566 -7 25612 273
rect 25824 -7 25870 273
rect 14622 -54 25870 -7
rect 14622 -55 14926 -54
rect 14622 -211 14668 -55
rect 14880 -211 14926 -55
rect 14622 -258 14926 -211
rect 14622 -539 14668 -258
rect 14880 -299 14926 -258
rect 14880 -499 15154 -299
rect 14880 -539 14926 -499
rect 14622 -586 14926 -539
rect 16580 -540 16976 -211
rect 18356 -499 18366 -299
rect 18418 -499 18428 -299
rect 18538 -500 18622 -54
rect 20120 -540 20516 -210
rect 21842 -499 21852 -299
rect 21904 -499 21914 -299
rect 22064 -499 22074 -299
rect 22126 -499 22136 -299
rect 23640 -540 24036 -210
rect 25566 -211 25612 -54
rect 25824 -211 25870 -54
rect 25566 -258 25870 -211
rect 25566 -299 25612 -258
rect 25338 -499 25612 -299
rect 25566 -539 25612 -499
rect 25824 -539 25870 -258
rect 14622 -743 14668 -586
rect 14880 -743 14926 -586
rect 14622 -790 14926 -743
rect 15164 -790 25328 -540
rect 25566 -586 25870 -539
rect 25566 -743 25612 -586
rect 25824 -743 25870 -586
rect 25566 -790 25870 -743
rect 14622 -1071 14668 -790
rect 14880 -831 14926 -790
rect 14880 -1031 15154 -831
rect 14880 -1071 14926 -1031
rect 14622 -1118 14926 -1071
rect 16580 -1118 16976 -790
rect 18356 -1031 18366 -830
rect 18418 -1031 18428 -830
rect 18578 -1031 18588 -831
rect 18640 -1031 18650 -831
rect 20120 -1118 20516 -790
rect 14622 -1276 14668 -1118
rect 14880 -1276 14926 -1118
rect 21870 -1276 21954 -830
rect 22064 -1031 22074 -831
rect 22126 -1031 22136 -831
rect 23641 -1118 24037 -790
rect 25566 -831 25612 -790
rect 25338 -1031 25612 -831
rect 25566 -1071 25612 -1031
rect 25824 -1071 25870 -790
rect 25566 -1118 25870 -1071
rect 25566 -1276 25612 -1118
rect 25824 -1276 25870 -1118
rect 14622 -1323 25870 -1276
rect 14622 -1603 14668 -1323
rect 14880 -1603 14926 -1323
rect 15108 -1602 15154 -1323
rect 15088 -1603 15154 -1602
rect 25566 -1603 25612 -1323
rect 25824 -1603 25870 -1323
rect 14622 -1649 25870 -1603
rect 14622 -1650 15088 -1649
rect 15134 -1650 25870 -1649
rect 16178 -2670 16224 -2637
rect 18089 -2670 18485 -2360
rect 20821 -2454 25839 -2408
rect 16178 -2778 20226 -2670
rect 16234 -2920 20226 -2778
rect 20821 -2718 20867 -2454
rect 21079 -2718 21125 -2454
rect 25535 -2718 25581 -2454
rect 25793 -2718 25839 -2454
rect 20821 -2764 25839 -2718
rect 18089 -3230 18485 -2920
rect 20821 -2994 20867 -2764
rect 21079 -2994 21125 -2764
rect 20821 -3040 20896 -2994
rect 21063 -3040 21125 -2994
rect 20821 -3364 20867 -3040
rect 21079 -3364 21125 -3040
rect 21443 -3332 21453 -3072
rect 21505 -3332 21515 -3072
rect 20821 -3410 20883 -3364
rect 21054 -3410 21125 -3364
rect 22118 -3410 22514 -2993
rect 23107 -3332 23117 -3072
rect 23169 -3332 23179 -3072
rect 23481 -3332 23491 -3072
rect 23543 -3332 23553 -3072
rect 20821 -3640 20867 -3410
rect 21079 -3640 21125 -3410
rect 22776 -3481 22963 -3410
rect 23615 -3413 23625 -3361
rect 23962 -3413 23972 -3361
rect 24262 -3410 24658 -2993
rect 25535 -2994 25581 -2764
rect 25793 -2994 25839 -2764
rect 25535 -3040 25605 -2994
rect 25769 -3040 25839 -2994
rect 25145 -3332 25155 -3072
rect 25207 -3332 25217 -3072
rect 25535 -3364 25581 -3040
rect 25793 -3364 25839 -3040
rect 25535 -3410 25601 -3364
rect 25770 -3410 25839 -3364
rect 22776 -3566 23882 -3481
rect 20821 -3686 20886 -3640
rect 21055 -3686 21125 -3640
rect 20821 -4010 20867 -3686
rect 21079 -4010 21125 -3686
rect 21443 -3978 21453 -3718
rect 21505 -3978 21515 -3718
rect 20821 -4056 20895 -4010
rect 21050 -4056 21125 -4010
rect 22113 -4056 22509 -3639
rect 22688 -3689 22698 -3637
rect 23035 -3689 23045 -3637
rect 23695 -3640 23882 -3566
rect 23107 -3978 23117 -3718
rect 23169 -3978 23179 -3718
rect 23481 -3978 23491 -3718
rect 23543 -3978 23553 -3718
rect 24262 -4056 24658 -3639
rect 25535 -3640 25581 -3410
rect 25793 -3640 25839 -3410
rect 25535 -3686 25599 -3640
rect 25767 -3686 25839 -3640
rect 25145 -3978 25155 -3718
rect 25207 -3978 25217 -3718
rect 25535 -4010 25581 -3686
rect 25793 -4010 25839 -3686
rect 25535 -4056 25607 -4010
rect 25765 -4056 25839 -4010
rect 20821 -4286 20867 -4056
rect 21079 -4286 21125 -4056
rect 25535 -4286 25581 -4056
rect 25793 -4286 25839 -4056
rect 20821 -4332 25839 -4286
rect 20821 -4596 20867 -4332
rect 21079 -4596 21125 -4332
rect 25535 -4596 25581 -4332
rect 25793 -4596 25839 -4332
rect 20821 -4642 25839 -4596
<< via1 >>
rect 21788 1989 21840 2189
rect 25338 1989 25390 2189
rect 21788 1458 21840 1657
rect 25338 1456 25390 1657
rect 18366 -499 18418 -299
rect 21852 -499 21904 -299
rect 22074 -499 22126 -299
rect 18366 -1031 18418 -830
rect 18588 -1031 18640 -831
rect 22074 -1031 22126 -831
rect 21453 -3332 21505 -3072
rect 23117 -3332 23169 -3072
rect 23491 -3332 23543 -3072
rect 23625 -3413 23962 -3361
rect 25155 -3332 25207 -3072
rect 21453 -3978 21505 -3718
rect 22698 -3689 23035 -3637
rect 23117 -3978 23169 -3718
rect 23491 -3978 23543 -3718
rect 25155 -3978 25207 -3718
<< metal2 >>
rect 21729 2388 25441 2398
rect 21896 2325 25274 2388
rect 21729 2315 25441 2325
rect 21786 2189 21842 2199
rect 21786 1979 21842 1989
rect 25338 2189 25390 2199
rect 25390 2042 26105 2052
rect 25390 1989 25525 2042
rect 25338 1979 25525 1989
rect 25692 1979 26105 2042
rect 25338 1969 26105 1979
rect 25585 1968 25645 1969
rect 21786 1657 21842 1667
rect 21786 1448 21842 1458
rect 25336 1657 25392 1667
rect 25336 1446 25392 1456
rect 21732 1327 21899 1337
rect 25515 1327 25682 1337
rect 21899 1263 25515 1327
rect 21732 1253 21899 1263
rect 25515 1253 25682 1263
rect 18309 575 22183 585
rect 18476 511 22016 575
rect 18309 501 22183 511
rect 18537 -104 26088 -94
rect 18704 -168 21791 -104
rect 21958 -168 26088 -104
rect 18537 -178 26088 -168
rect 25898 -179 26088 -178
rect 18364 -299 18420 -289
rect 18364 -509 18420 -499
rect 21850 -299 21906 -289
rect 21850 -509 21906 -499
rect 22072 -299 22128 -289
rect 22072 -509 22128 -499
rect 18364 -830 18420 -820
rect 18364 -1041 18420 -1031
rect 18586 -831 18642 -821
rect 18586 -1041 18642 -1031
rect 22072 -831 22128 -821
rect 22072 -1042 22128 -1032
rect 26061 -2807 26125 -2797
rect 21397 -2847 26061 -2837
rect 21564 -2911 26061 -2847
rect 21397 -2921 26061 -2911
rect 26061 -2984 26125 -2974
rect 21451 -3072 21507 -3062
rect 21451 -3342 21507 -3332
rect 23115 -3072 23171 -3062
rect 23115 -3342 23171 -3332
rect 23489 -3072 23545 -3062
rect 23489 -3342 23545 -3332
rect 25153 -3072 25209 -3062
rect 25153 -3343 25209 -3333
rect 23625 -3359 23962 -3349
rect 23625 -3425 23962 -3415
rect 22786 -3483 23775 -3482
rect 22786 -3492 23872 -3483
rect 22953 -3493 23872 -3492
rect 22953 -3556 23705 -3493
rect 22786 -3557 23705 -3556
rect 22786 -3566 23872 -3557
rect 23705 -3567 23872 -3566
rect 22698 -3635 23035 -3625
rect 22698 -3701 23035 -3691
rect 21451 -3718 21507 -3708
rect 21451 -3988 21507 -3978
rect 23115 -3718 23171 -3708
rect 23115 -3988 23171 -3978
rect 23489 -3718 23545 -3708
rect 23489 -3988 23545 -3978
rect 25155 -3718 25207 -3708
rect 26061 -3771 26125 -3761
rect 25207 -3889 26061 -3805
rect 26061 -3948 26125 -3938
rect 25155 -3988 25207 -3978
rect 21422 -4139 25259 -4129
rect 21422 -4203 21428 -4139
rect 21595 -4203 25092 -4139
rect 21422 -4213 25259 -4203
<< via2 >>
rect 21729 2325 21896 2388
rect 25274 2325 25441 2388
rect 21786 1989 21788 2189
rect 21788 1989 21840 2189
rect 21840 1989 21842 2189
rect 25525 1979 25692 2042
rect 21786 1458 21788 1657
rect 21788 1458 21840 1657
rect 21840 1458 21842 1657
rect 25336 1456 25338 1657
rect 25338 1456 25390 1657
rect 25390 1456 25392 1657
rect 21732 1263 21899 1327
rect 25515 1263 25682 1327
rect 18309 511 18476 575
rect 22016 511 22183 575
rect 18537 -168 18704 -104
rect 21791 -168 21958 -104
rect 18364 -499 18366 -299
rect 18366 -499 18418 -299
rect 18418 -499 18420 -299
rect 21850 -499 21852 -299
rect 21852 -499 21904 -299
rect 21904 -499 21906 -299
rect 22072 -499 22074 -299
rect 22074 -499 22126 -299
rect 22126 -499 22128 -299
rect 18364 -1031 18366 -830
rect 18366 -1031 18418 -830
rect 18418 -1031 18420 -830
rect 18586 -1031 18588 -831
rect 18588 -1031 18640 -831
rect 18640 -1031 18642 -831
rect 22072 -1031 22074 -831
rect 22074 -1031 22126 -831
rect 22126 -1031 22128 -831
rect 22072 -1032 22128 -1031
rect 21397 -2911 21564 -2847
rect 26061 -2974 26125 -2807
rect 21451 -3332 21453 -3072
rect 21453 -3332 21505 -3072
rect 21505 -3332 21507 -3072
rect 23115 -3332 23117 -3072
rect 23117 -3332 23169 -3072
rect 23169 -3332 23171 -3072
rect 23489 -3332 23491 -3072
rect 23491 -3332 23543 -3072
rect 23543 -3332 23545 -3072
rect 25153 -3332 25155 -3072
rect 25155 -3332 25207 -3072
rect 25207 -3332 25209 -3072
rect 25153 -3333 25209 -3332
rect 23625 -3361 23962 -3359
rect 23625 -3413 23962 -3361
rect 23625 -3415 23962 -3413
rect 22786 -3556 22953 -3492
rect 23705 -3557 23872 -3493
rect 22698 -3637 23035 -3635
rect 22698 -3689 23035 -3637
rect 22698 -3691 23035 -3689
rect 21451 -3978 21453 -3718
rect 21453 -3978 21505 -3718
rect 21505 -3978 21507 -3718
rect 23115 -3978 23117 -3718
rect 23117 -3978 23169 -3718
rect 23169 -3978 23171 -3718
rect 23489 -3978 23491 -3718
rect 23491 -3978 23543 -3718
rect 23543 -3978 23545 -3718
rect 26061 -3938 26125 -3771
rect 21428 -4203 21595 -4139
rect 25092 -4203 25259 -4139
<< metal3 >>
rect 21719 2388 21906 2393
rect 21719 2325 21729 2388
rect 21896 2325 21906 2388
rect 21719 2320 21906 2325
rect 25264 2388 25451 2393
rect 25264 2325 25274 2388
rect 25441 2325 25451 2388
rect 25264 2320 25451 2325
rect 21776 2189 21852 2320
rect 21776 1989 21786 2189
rect 21842 1989 21852 2189
rect 21776 1984 21852 1989
rect 21776 1657 21852 1662
rect 21776 1458 21786 1657
rect 21842 1458 21852 1657
rect 21776 1332 21852 1458
rect 25326 1657 25402 2320
rect 25515 2042 25702 2047
rect 25515 1979 25525 2042
rect 25692 1979 25702 2042
rect 25515 1974 25702 1979
rect 25326 1456 25336 1657
rect 25392 1456 25402 1657
rect 25326 1451 25402 1456
rect 25583 1332 25647 1974
rect 21722 1327 21909 1332
rect 21722 1263 21732 1327
rect 21899 1263 21909 1327
rect 21722 1258 21909 1263
rect 25505 1327 25692 1332
rect 25505 1263 25515 1327
rect 25682 1263 25692 1327
rect 25505 1258 25692 1263
rect 18299 575 18486 580
rect 18299 511 18309 575
rect 18476 511 18486 575
rect 18299 506 18486 511
rect 22006 575 22193 580
rect 22006 511 22016 575
rect 22183 511 22193 575
rect 22006 506 22193 511
rect 18354 -299 18430 506
rect 18527 -104 18714 -99
rect 18527 -168 18537 -104
rect 18704 -168 18714 -104
rect 18527 -173 18714 -168
rect 21781 -104 21968 -99
rect 21781 -168 21791 -104
rect 21958 -168 21968 -104
rect 21781 -173 21968 -168
rect 18354 -499 18364 -299
rect 18420 -499 18430 -299
rect 18354 -830 18430 -499
rect 18354 -1031 18364 -830
rect 18420 -1031 18430 -830
rect 18354 -1036 18430 -1031
rect 18576 -831 18652 -173
rect 21840 -299 21916 -173
rect 21840 -499 21850 -299
rect 21906 -499 21916 -299
rect 21840 -504 21916 -499
rect 22062 -299 22138 506
rect 22062 -499 22072 -299
rect 22128 -499 22138 -299
rect 18576 -1031 18586 -831
rect 18642 -1031 18652 -831
rect 18576 -1036 18652 -1031
rect 22062 -831 22138 -499
rect 22062 -1032 22072 -831
rect 22128 -1032 22138 -831
rect 22062 -1037 22138 -1032
rect 26051 -2807 26135 -2802
rect 21387 -2847 21574 -2842
rect 21387 -2911 21397 -2847
rect 21564 -2911 21574 -2847
rect 21387 -2916 21574 -2911
rect 21441 -3072 21517 -2916
rect 26051 -2974 26061 -2807
rect 26125 -2974 26135 -2807
rect 21441 -3332 21451 -3072
rect 21507 -3332 21517 -3072
rect 21441 -3337 21517 -3332
rect 23105 -3072 23555 -3067
rect 23105 -3332 23115 -3072
rect 23171 -3332 23489 -3072
rect 23545 -3332 23555 -3072
rect 22776 -3492 22963 -3487
rect 22776 -3556 22786 -3492
rect 22953 -3556 22963 -3492
rect 22776 -3630 22963 -3556
rect 22688 -3635 23045 -3630
rect 22688 -3691 22698 -3635
rect 23035 -3691 23045 -3635
rect 22688 -3696 23045 -3691
rect 21441 -3718 21517 -3713
rect 21441 -3978 21451 -3718
rect 21507 -3978 21517 -3718
rect 21441 -4134 21517 -3978
rect 23105 -3718 23555 -3332
rect 25143 -3072 25219 -3067
rect 25143 -3333 25153 -3072
rect 25209 -3333 25219 -3072
rect 23615 -3359 23972 -3354
rect 23615 -3415 23625 -3359
rect 23962 -3415 23972 -3359
rect 23615 -3420 23972 -3415
rect 23695 -3493 23882 -3420
rect 23695 -3557 23705 -3493
rect 23872 -3557 23882 -3493
rect 23695 -3562 23882 -3557
rect 23105 -3978 23115 -3718
rect 23171 -3978 23489 -3718
rect 23545 -3978 23555 -3718
rect 23105 -3983 23555 -3978
rect 25143 -4134 25219 -3333
rect 26051 -3771 26135 -2974
rect 26051 -3938 26061 -3771
rect 26125 -3938 26135 -3771
rect 26051 -3943 26135 -3938
rect 21418 -4139 21605 -4134
rect 21418 -4203 21428 -4139
rect 21595 -4203 21605 -4139
rect 21418 -4208 21605 -4203
rect 25082 -4139 25269 -4134
rect 25082 -4203 25092 -4139
rect 25259 -4203 25269 -4139
rect 25082 -4208 25269 -4203
use trans_gate  x1
timestamp 1711994542
transform 1 0 11684 0 1 -1512
box 0 -2380 2272 590
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[0]
timestamp 1712074089
transform 1 0 21460 0 1 2621
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[1]
timestamp 1712074089
transform 1 0 21460 0 1 2089
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[2]
timestamp 1712074089
transform 1 0 21460 0 1 1557
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XDM1[3]
timestamp 1712074089
transform 1 0 21460 0 1 1025
box -296 -319 296 319
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[0]
timestamp 1712318662
transform 1 0 24349 0 1 -3848
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM1[1]
timestamp 1712318662
transform 1 0 22311 0 1 -3202
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM2[0]
timestamp 1712318662
transform 1 0 24349 0 1 -3202
box -1028 -388 1028 388
use sky130_fd_pr__nfet_g5v0d10v5_LQ7VVE  XM2[1]
timestamp 1712318662
transform 1 0 22311 0 1 -3848
box -1028 -388 1028 388
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[0]
timestamp 1712064068
transform -1 0 22646 0 -1 1557
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM3[1]
timestamp 1712064068
transform 1 0 24532 0 1 2089
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[0]
timestamp 1712319635
transform 1 0 20246 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM4[1]
timestamp 1712319635
transform 1 0 20246 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[0]
timestamp 1712064068
transform 1 0 24532 0 1 1557
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XM5[1]
timestamp 1712064068
transform 1 0 22646 0 1 2089
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[0]
timestamp 1712319635
transform 1 0 16760 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[1]
timestamp 1712319635
transform 1 0 16760 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[2]
timestamp 1712319635
transform 1 0 23732 0 1 -399
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XM6[3]
timestamp 1712319635
transform 1 0 23732 0 1 -931
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_GGMWVD  XM7
timestamp 1711994542
transform 0 1 26587 -1 0 1944
box -996 -319 996 319
use sky130_fd_pr__nfet_01v8_L8NDKD  XM8
timestamp 1712242108
transform 0 1 26578 -1 0 -2708
box -996 -310 996 310
use sky130_fd_pr__pfet_01v8_3HBZVM  XM9
timestamp 1711994542
transform 1 0 26564 0 1 175
box -296 -519 296 519
use sky130_fd_pr__nfet_01v8_C8TQ3N  XM10
timestamp 1711994542
transform 1 0 26564 0 1 -1094
box -296 -510 296 510
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM11
timestamp 1712318662
transform 1 0 18230 0 1 -2538
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_7ZF23Z  XM12
timestamp 1712318662
transform 1 0 18230 0 1 -3052
box -2196 -310 2196 310
use sky130_fd_pr__nfet_01v8_V433WY  XM13
timestamp 1711994542
transform -1 0 19928 0 -1 -3997
box -496 -310 496 310
use sky130_fd_pr__nfet_01v8_V433WY  XM14
timestamp 1711994542
transform -1 0 19928 0 -1 -4511
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM15
timestamp 1711994542
transform 1 0 20414 0 1 1025
box -496 -319 496 319
use sky130_fd_pr__pfet_01v8_C2YSV5  XM16
timestamp 1711994542
transform 1 0 20414 0 1 1557
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM17
timestamp 1711994542
transform 0 1 26578 -1 0 -4326
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_C2YSV5  XM18
timestamp 1711994542
transform 1 0 14974 0 1 -2547
box -496 -319 496 319
use sky130_fd_pr__nfet_01v8_V433WY  XM19
timestamp 1711994542
transform 1 0 14988 0 1 -3282
box -496 -310 496 310
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[4]
timestamp 1712074089
transform 1 0 25718 0 1 2621
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[5]
timestamp 1712074089
transform 1 0 25718 0 1 2089
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[6]
timestamp 1712074089
transform 1 0 25718 0 1 1557
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[7]
timestamp 1712074089
transform 1 0 25718 0 1 1025
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[8]
timestamp 1712074089
transform 1 0 14774 0 1 133
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[9]
timestamp 1712074089
transform 1 0 14774 0 1 -399
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[10]
timestamp 1712074089
transform 1 0 14774 0 1 -931
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[11]
timestamp 1712074089
transform 1 0 14774 0 1 -1463
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[12]
timestamp 1712074089
transform 1 0 25718 0 1 133
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[13]
timestamp 1712074089
transform 1 0 25718 0 1 -399
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[14]
timestamp 1712074089
transform 1 0 25718 0 1 -931
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_J2L9E5  XMD1[15]
timestamp 1712074089
transform 1 0 25718 0 1 -1463
box -296 -319 296 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[0]
timestamp 1712319635
transform 1 0 16760 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[1]
timestamp 1712319635
transform 1 0 20246 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[2]
timestamp 1712319635
transform 1 0 23732 0 1 133
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[3]
timestamp 1712319635
transform 1 0 16760 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[4]
timestamp 1712319635
transform 1 0 20246 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_XTWSDC  XMD16[5]
timestamp 1712319635
transform 1 0 23732 0 1 -1463
box -1796 -319 1796 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[0]
timestamp 1712064068
transform 1 0 22646 0 1 2621
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[1]
timestamp 1712064068
transform 1 0 24532 0 1 2621
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[2]
timestamp 1712064068
transform 1 0 22646 0 1 1025
box -996 -319 996 319
use sky130_fd_pr__pfet_01v8_G3L97A  XMD[3]
timestamp 1712064068
transform 1 0 24532 0 1 1025
box -996 -319 996 319
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[0]
timestamp 1712318662
transform 1 0 20973 0 1 -2586
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[1]
timestamp 1712318662
transform 1 0 20973 0 1 -4464
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[2]
timestamp 1712318662
transform 1 0 25687 0 1 -2586
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_CD9S2Z  XMDN1[3]
timestamp 1712318662
transform 1 0 25687 0 1 -4464
box -328 -358 328 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[0]
timestamp 1712318662
transform 1 0 22311 0 1 -2586
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[1]
timestamp 1712318662
transform 1 0 24349 0 1 -2586
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[2]
timestamp 1712318662
transform 1 0 22311 0 1 -4464
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_DEN7YK  XMDN8[3]
timestamp 1712318662
transform 1 0 24349 0 1 -4464
box -1028 -358 1028 358
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[0]
timestamp 1712318662
transform 1 0 20973 0 1 -3202
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[1]
timestamp 1712318662
transform 1 0 20973 0 1 -3848
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[2]
timestamp 1712318662
transform 1 0 25687 0 1 -3202
box -328 -388 328 388
use sky130_fd_pr__nfet_g5v0d10v5_4T6WVE  XMDN13[3]
timestamp 1712318662
transform 1 0 25687 0 1 -3848
box -328 -388 328 388
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1713529122
<< dnwell >>
rect -18138 9035 5931 17409
rect 7922 10297 23998 15120
rect -18138 -3922 10182 9035
rect 11442 -336 23998 10297
<< nwell >>
rect -18218 17203 6011 17489
rect -18218 -3716 -17932 17203
rect 5725 9115 6011 17203
rect 7842 14914 24078 15200
rect 7842 10503 8128 14914
rect 7842 10217 11648 10503
rect 5725 8829 10262 9115
rect 9976 -3716 10262 8829
rect 11362 -130 11648 10217
rect 23792 -130 24078 14914
rect 11362 -416 24078 -130
rect -18218 -4002 10262 -3716
<< nsubdiff >>
rect -18182 17433 5975 17453
rect -18182 17399 -18100 17433
rect 5895 17399 5975 17433
rect -18182 17379 5975 17399
rect -18182 17373 -18108 17379
rect -18182 -3883 -18162 17373
rect -18128 -3883 -18108 17373
rect 5901 17375 5975 17379
rect 5901 9087 5921 17375
rect 5955 9087 5975 17375
rect 7878 15144 24042 15164
rect 7878 15110 8003 15144
rect 23965 15110 24042 15144
rect 7878 15090 24042 15110
rect 7878 15084 8001 15090
rect 7878 10333 7898 15084
rect 7932 10333 8001 15084
rect 7878 10327 8001 10333
rect 23968 15084 24042 15090
rect 7878 10307 11473 10327
rect 7878 10273 8004 10307
rect 11397 10273 11473 10307
rect 7878 10253 11473 10273
rect 5901 9079 5975 9087
rect 11399 10247 11473 10253
rect 5901 9059 10225 9079
rect 5901 9025 5976 9059
rect 10148 9025 10225 9059
rect 5901 9005 10225 9025
rect -18182 -3891 -18108 -3883
rect 10151 8999 10225 9005
rect 10151 -3885 10171 8999
rect 10205 -3885 10225 8999
rect 11399 -299 11419 10247
rect 11453 -299 11473 10247
rect 11399 -305 11473 -299
rect 23968 -297 23988 15084
rect 24022 -297 24042 15084
rect 23968 -305 24042 -297
rect 11399 -325 24042 -305
rect 11399 -359 11479 -325
rect 23968 -359 24042 -325
rect 11399 -379 24042 -359
rect 10151 -3891 10225 -3885
rect -18182 -3912 10225 -3891
rect -18182 -3946 -18108 -3912
rect 10145 -3946 10225 -3912
rect -18182 -3966 10225 -3946
<< nsubdiffcont >>
rect -18100 17399 5895 17433
rect -18162 -3883 -18128 17373
rect 5921 9087 5955 17375
rect 8003 15110 23965 15144
rect 7898 10333 7932 15084
rect 8004 10273 11397 10307
rect 5976 9025 10148 9059
rect 10171 -3885 10205 8999
rect 11419 -299 11453 10247
rect 23988 -297 24022 15084
rect 11479 -359 23968 -325
rect -18108 -3946 10145 -3912
<< locali >>
rect -18162 17399 -18100 17433
rect 5895 17399 5955 17433
rect -18162 17373 -18128 17399
rect 5921 17375 5955 17399
rect 7898 15110 8003 15144
rect 23965 15110 24022 15144
rect 7898 15084 7932 15110
rect 7898 10307 7932 10333
rect 23988 15084 24022 15110
rect 7898 10273 8004 10307
rect 11397 10273 11453 10307
rect 5921 9059 5955 9087
rect 11419 10247 11453 10273
rect 5921 9025 5976 9059
rect 10148 9025 10205 9059
rect -18162 -3912 -18128 -3883
rect 10171 8999 10205 9025
rect 13561 6483 15409 6488
rect 11419 -325 11453 -299
rect 23988 -325 24022 -297
rect 11419 -359 11479 -325
rect 23968 -359 24022 -325
rect 10171 -3912 10205 -3885
rect -18162 -3946 -18108 -3912
rect 10145 -3946 10205 -3912
<< metal1 >>
rect -18218 16076 5440 17489
rect 7535 17445 24079 17489
rect -17312 16075 5440 16076
rect 7380 16078 24079 17445
rect -1954 13119 -1838 16075
rect -320 13119 -204 16075
rect 1358 13119 1474 16075
rect 3026 11509 3142 16075
rect -448 9664 -438 9804
rect -381 9664 -371 9804
rect 1230 8849 1240 8989
rect 1297 8849 1307 8989
rect 4779 8827 4977 16075
rect 7380 15179 7927 16078
rect 7380 10253 7878 15179
rect 13852 13450 16007 16078
rect 23199 10475 23247 10653
rect 7380 9756 11694 10253
rect 7380 9746 7877 9756
rect 4779 8629 7597 8827
rect 7399 8476 7597 8629
rect 11104 8476 11694 9756
rect 7399 8277 7722 8476
rect 11104 8278 11976 8476
rect 7399 6284 7597 8277
rect 9759 6502 10025 6701
rect 7399 6085 7723 6284
rect 2897 4025 2907 4165
rect 2964 4025 2974 4165
rect -854 -2701 -738 299
rect 780 -2701 896 299
rect 2458 -2701 2574 299
rect 4126 -2701 4242 1909
rect 4547 1590 4685 4904
rect 7399 4092 7597 6085
rect 9826 4509 10025 6502
rect 9759 4310 10025 4509
rect 7399 3894 7775 4092
rect 7399 1900 7597 3894
rect 9826 2317 10025 4310
rect 9759 2118 10025 2317
rect 7399 1701 7702 1900
rect 4535 1533 4545 1590
rect 4685 1533 4695 1590
rect 9826 125 10025 2118
rect 11104 6284 11694 8278
rect 13706 7672 13824 7682
rect 13706 7616 13717 7672
rect 13857 7616 13867 7672
rect 13706 7606 13824 7616
rect 13706 7605 13857 7606
rect 12737 6502 13315 6782
rect 13035 6487 13315 6502
rect 11104 6086 11966 6284
rect 13035 6207 13316 6487
rect 11104 4092 11694 6086
rect 13035 4589 13315 6207
rect 11753 4310 13315 4589
rect 11104 3894 11965 4092
rect 11104 1900 11694 3894
rect 13035 2397 13315 4310
rect 11753 2118 13315 2397
rect 11104 1702 11946 1900
rect 13035 206 13315 2118
rect 9759 -74 10025 125
rect 11753 -73 13315 206
rect 9826 -2701 10025 -74
rect 13035 -2700 13315 -73
rect 15779 -2700 17934 6277
rect -18218 -4002 10025 -2701
rect 13032 -2705 17934 -2700
rect 13032 -4002 24405 -2705
<< via1 >>
rect -438 9664 -381 9804
rect 1240 8849 1297 8989
rect 22900 10492 23196 10635
rect 5953 6328 6147 6436
rect 2907 4025 2964 4165
rect 4545 1533 4685 1590
rect 13717 7616 13857 7672
<< metal2 >>
rect 22876 10635 24078 10653
rect 22876 10492 22900 10635
rect 23196 10492 24078 10635
rect 22876 10475 24078 10492
rect 7296 10417 13114 10422
rect 7296 10414 12960 10417
rect 7296 10358 7308 10414
rect 7448 10361 12960 10414
rect 13100 10361 13114 10417
rect 7448 10358 13114 10361
rect 7296 10348 13114 10358
rect -438 9804 -381 9814
rect -381 9765 7502 9775
rect -381 9708 7362 9765
rect -381 9698 7502 9708
rect -438 9654 -381 9664
rect -438 9337 -381 9347
rect -381 9298 7292 9308
rect -381 9241 7142 9298
rect 7282 9241 7292 9298
rect -381 9231 7292 9241
rect -438 9187 -381 9197
rect 1240 8989 1297 8999
rect 1297 8951 7071 8961
rect 1297 8894 6920 8951
rect 7060 8894 7071 8951
rect 1297 8884 7071 8894
rect 1240 8839 1297 8849
rect 1240 8541 1297 8551
rect 1230 8433 1240 8510
rect 1297 8500 6847 8510
rect 1297 8443 6697 8500
rect 6837 8443 6847 8500
rect 1297 8433 6847 8443
rect 1240 8391 1297 8401
rect 7352 8170 7882 8173
rect 7352 8163 7892 8170
rect 7352 8106 7362 8163
rect 7502 8106 7892 8163
rect 7352 8099 7892 8106
rect 7352 8096 7882 8099
rect 12950 7672 13857 7682
rect 12950 7616 12962 7672
rect 13102 7616 13717 7672
rect 12950 7605 13857 7616
rect 7131 7563 7882 7569
rect 7131 7556 7934 7563
rect 7131 7499 7142 7556
rect 7282 7499 7934 7556
rect 7131 7497 7934 7499
rect 7131 7492 7882 7497
rect 13261 7203 13669 7207
rect 13261 7189 13672 7203
rect 13261 7081 13268 7189
rect 13462 7081 13672 7189
rect 13261 7054 13672 7081
rect 13261 7047 13669 7054
rect 11196 6968 11894 6978
rect 11196 6890 11209 6968
rect 11349 6890 11894 6968
rect 11196 6880 11894 6890
rect 5947 6436 13159 6442
rect 5947 6328 5953 6436
rect 6147 6328 12956 6436
rect 13150 6328 13159 6436
rect 5947 6322 13159 6328
rect 12951 6106 23104 6111
rect 12951 5998 12960 6106
rect 13154 6097 23104 6106
rect 13154 6006 22940 6097
rect 23093 6006 23104 6097
rect 13154 5998 23104 6006
rect 12951 5991 23104 5998
rect 6910 5974 7882 5981
rect 6910 5971 7903 5974
rect 6910 5914 6920 5971
rect 7060 5914 7903 5971
rect 6910 5904 7903 5914
rect 20888 5941 23283 5942
rect 20888 5928 24078 5941
rect 20888 5837 20901 5928
rect 21054 5837 24078 5928
rect 20888 5822 24078 5837
rect 23283 5821 24078 5822
rect 6686 5372 7882 5377
rect 6686 5367 7969 5372
rect 6686 5310 6697 5367
rect 6837 5310 7969 5367
rect 6686 5305 7969 5310
rect 6686 5300 7882 5305
rect 10860 4776 11911 4786
rect 10860 4698 10873 4776
rect 11013 4698 11911 4776
rect 10860 4688 11911 4698
rect 2907 4165 2964 4175
rect 2964 4131 7362 4142
rect 2964 4121 7512 4131
rect 2964 4065 7362 4121
rect 7502 4064 7512 4121
rect 7362 4054 7512 4064
rect 2907 4015 2964 4025
rect 7352 3783 7882 3789
rect 7352 3779 7939 3783
rect 2907 3713 2964 3723
rect 7352 3722 7362 3779
rect 7502 3722 7939 3779
rect 7352 3721 7939 3722
rect 7352 3713 7882 3721
rect 7362 3712 7502 3713
rect 7576 3712 7882 3713
rect 2964 3670 7292 3680
rect 2964 3613 7142 3670
rect 7282 3613 7292 3670
rect 2964 3603 7292 3613
rect 2907 3563 2964 3573
rect 7132 3181 7882 3185
rect 7132 3175 7903 3181
rect 7132 3118 7142 3175
rect 7282 3118 7903 3175
rect 7132 3108 7903 3118
rect 10555 2584 11866 2594
rect 10555 2506 10568 2584
rect 10708 2506 11866 2584
rect 10555 2496 11866 2506
rect 4537 1597 4674 1600
rect 4537 1590 7886 1597
rect 4537 1533 4545 1590
rect 4685 1533 7919 1590
rect 4537 1527 7919 1533
rect 4537 1523 7886 1527
rect 4537 636 7882 638
rect 4537 629 7898 636
rect 4537 572 4546 629
rect 4686 597 7898 629
rect 4686 572 8482 597
rect 4537 566 8482 572
rect 10263 392 11995 402
rect 10263 314 10276 392
rect 10416 314 11995 392
rect 10263 304 11995 314
rect -2050 -1881 13469 -1859
rect -2050 -2046 13294 -1881
rect 13434 -2046 13469 -1881
rect -2050 -2079 13469 -2046
<< via2 >>
rect 7308 10358 7448 10414
rect 12960 10361 13100 10417
rect 7362 9708 7502 9765
rect -438 9197 -381 9337
rect 7142 9241 7282 9298
rect 6920 8894 7060 8951
rect 1240 8401 1297 8541
rect 6697 8443 6837 8500
rect 7362 8106 7502 8163
rect 12962 7616 13102 7672
rect 7142 7499 7282 7556
rect 13268 7081 13462 7189
rect 11209 6890 11349 6968
rect 12956 6328 13150 6436
rect 12960 5998 13154 6106
rect 22940 6006 23093 6097
rect 6920 5914 7060 5971
rect 20901 5837 21054 5928
rect 6697 5310 6837 5367
rect 10873 4698 11013 4776
rect 7362 4064 7502 4121
rect 7362 3722 7502 3779
rect 2907 3573 2964 3713
rect 7142 3613 7282 3670
rect 7142 3118 7282 3175
rect 10568 2506 10708 2584
rect 4546 572 4686 629
rect 10276 314 10416 392
rect 13294 -2046 13434 -1881
<< metal3 >>
rect 7296 10414 7460 17924
rect 7296 10358 7308 10414
rect 7448 10358 7460 10414
rect 7296 10348 7460 10358
rect 12950 10417 13114 10422
rect 12950 10361 12960 10417
rect 13100 10361 13114 10417
rect 7352 9765 7512 9775
rect 7352 9708 7362 9765
rect 7502 9708 7512 9765
rect -448 9337 -371 9342
rect -448 9197 -438 9337
rect -381 9197 -371 9337
rect -448 9192 -371 9197
rect 7131 9298 7292 9308
rect 7131 9241 7142 9298
rect 7282 9241 7292 9298
rect 6910 8951 7071 8961
rect 6910 8894 6920 8951
rect 7060 8894 7071 8951
rect 1230 8541 1307 8546
rect 1230 8401 1240 8541
rect 1297 8401 1307 8541
rect 1230 8396 1307 8401
rect 6686 8500 6847 8510
rect 6686 8443 6697 8500
rect 6837 8443 6847 8500
rect 6686 5367 6847 8443
rect 6910 5971 7071 8894
rect 7131 7556 7292 9241
rect 7352 8163 7512 9708
rect 7352 8106 7362 8163
rect 7502 8106 7512 8163
rect 7352 8096 7512 8106
rect 12950 7672 13114 10361
rect 12950 7616 12962 7672
rect 13102 7616 13114 7672
rect 12950 7605 13114 7616
rect 7131 7499 7142 7556
rect 7282 7499 7292 7556
rect 7131 7492 7292 7499
rect 13261 7189 13469 7207
rect 13261 7081 13268 7189
rect 13462 7081 13469 7189
rect 6910 5914 6920 5971
rect 7060 5914 7071 5971
rect 6910 5904 7071 5914
rect 11196 6968 11362 6978
rect 11196 6890 11209 6968
rect 11349 6890 11362 6968
rect 6686 5310 6697 5367
rect 6837 5310 6847 5367
rect 6686 5300 6847 5310
rect 4537 4901 4685 4974
rect 2897 3713 2974 3718
rect 2897 3573 2907 3713
rect 2964 3573 2974 3713
rect 2897 3568 2974 3573
rect 4537 629 4691 4901
rect 10860 4776 11026 4786
rect 10860 4698 10873 4776
rect 11013 4698 11026 4776
rect 7352 4121 7512 4131
rect 7352 4064 7362 4121
rect 7502 4064 7512 4121
rect 7352 3779 7512 4064
rect 7352 3722 7362 3779
rect 7502 3722 7512 3779
rect 7352 3713 7512 3722
rect 7132 3670 7292 3680
rect 7132 3613 7142 3670
rect 7282 3613 7292 3670
rect 7132 3175 7292 3613
rect 7132 3118 7142 3175
rect 7282 3118 7292 3175
rect 7132 3108 7292 3118
rect 4537 572 4546 629
rect 4686 572 4691 629
rect 4537 566 4691 572
rect 10555 2584 10721 2594
rect 10555 2506 10568 2584
rect 10708 2506 10721 2584
rect 10263 392 10429 402
rect 10263 314 10276 392
rect 10416 314 10429 392
rect 10263 -4002 10429 314
rect 10555 -4002 10721 2506
rect 10860 -4002 11026 4698
rect 11196 -420 11362 6890
rect 12951 6436 13159 6442
rect 12951 6328 12956 6436
rect 13150 6328 13159 6436
rect 12951 6106 13159 6328
rect 12951 5998 12960 6106
rect 13154 5998 13159 6106
rect 12951 5991 13159 5998
rect 11195 -4002 11361 -420
rect 13261 -1881 13469 7081
rect 20889 5928 21066 6265
rect 22927 6097 23104 6264
rect 22927 6006 22940 6097
rect 23093 6006 23104 6097
rect 22927 5991 23104 6006
rect 20889 5837 20901 5928
rect 21054 5837 21066 5928
rect 20889 5821 21066 5837
rect 13261 -2046 13294 -1881
rect 13434 -2046 13469 -1881
rect 13261 -4002 13469 -2046
<< fillblock >>
rect 18268 2356 20844 5659
rect 21598 101 23454 3000
use comp_hyst  comp_hyst_0
timestamp 1713226135
transform 1 0 6715 0 1 11492
box 1667 -5363 16947 2564
use initials  initials_0
timestamp 1713221383
transform 1 0 16849 0 1 2277
box 1419 79 3995 3382
use level_shifter  level_shifter_0
timestamp 1713359379
transform 1 0 6519 0 1 8816
box 1105 -2399 6458 -251
use level_shifter  level_shifter_1
timestamp 1713359379
transform 1 0 6519 0 1 6624
box 1105 -2399 6458 -251
use level_shifter  level_shifter_2
timestamp 1713359379
transform 1 0 6519 0 1 4432
box 1105 -2399 6458 -251
use level_shifter  level_shifter_3
timestamp 1713359379
transform 1 0 6519 0 1 2240
box 1105 -2399 6458 -251
use multiplexer  multiplexer_0
timestamp 1713226135
transform 1 0 -1955 0 1 209
box -199 -135 8108 13095
use rocket  rocket_0
timestamp 1713228654
transform 1 0 21607 0 1 457
box -9 -356 1847 2543
use vd2mux_conn  vd2mux_conn_1
timestamp 1713221383
transform 1 0 478 0 1 1
box -3578 973 -2488 12383
use voltage_divider  voltage_divider_0
timestamp 1713226135
transform 1 0 -16053 0 1 -2158
box -1259 -1438 14153 19128
<< labels >>
flabel metal3 7296 17760 7460 17924 0 FreeSans 1600 0 0 0 ibias
port 12 nsew
flabel metal2 13425 5991 22940 6111 0 FreeSans 800 0 0 0 vin
flabel metal1 -18218 -4002 10025 -2701 0 FreeSans 8000 0 0 0 avss
port 18 nsew
flabel metal1 -18218 16076 5440 17489 0 FreeSans 8000 0 0 0 avdd
port 15 nsew
flabel metal1 13032 -4002 24405 -2705 0 FreeSans 8000 0 0 0 dvss
port 16 nsew
flabel metal1 7535 16078 24079 17489 0 FreeSans 8000 0 0 0 dvdd
port 19 nsew
flabel metal3 10263 -4002 10429 -3847 0 FreeSans 1600 90 0 0 vtrip[3]
port 2 nsew
flabel metal3 10555 -4002 10721 -3848 0 FreeSans 1600 90 0 0 vtrip[2]
port 3 nsew
flabel metal3 10860 -4002 11026 -3848 0 FreeSans 1600 90 0 0 vtrip[1]
port 4 nsew
flabel metal3 11195 -4002 11361 -3848 0 FreeSans 1600 90 0 0 vtrip[0]
port 5 nsew
flabel metal3 13261 -4002 13469 -3848 0 FreeSans 1600 0 0 0 ena
port 17 nsew
flabel metal2 23788 5821 24078 5941 0 FreeSans 1600 0 0 0 vbg
port 10 nsew
flabel metal2 23196 10475 24078 10653 0 FreeSans 1600 0 0 0 ovout
port 20 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1712629466
<< xpolycontact >>
rect -9024 5150 -8742 5582
rect -9024 1930 -8742 2362
rect -8646 5150 -8364 5582
rect -8646 1930 -8364 2362
rect -8268 5150 -7986 5582
rect -8268 1930 -7986 2362
rect -7890 5150 -7608 5582
rect -7890 1930 -7608 2362
rect -7512 5150 -7230 5582
rect -7512 1930 -7230 2362
rect -7134 5150 -6852 5582
rect -7134 1930 -6852 2362
rect -6756 5150 -6474 5582
rect -6756 1930 -6474 2362
rect -6378 5150 -6096 5582
rect -6378 1930 -6096 2362
rect -6000 5150 -5718 5582
rect -6000 1930 -5718 2362
rect -5622 5150 -5340 5582
rect -5622 1930 -5340 2362
rect -5244 5150 -4962 5582
rect -5244 1930 -4962 2362
rect -4866 5150 -4584 5582
rect -4866 1930 -4584 2362
rect -4488 5150 -4206 5582
rect -4488 1930 -4206 2362
rect -4110 5150 -3828 5582
rect -4110 1930 -3828 2362
rect -3732 5150 -3450 5582
rect -3732 1930 -3450 2362
rect -3354 5150 -3072 5582
rect -3354 1930 -3072 2362
rect -2976 5150 -2694 5582
rect -2976 1930 -2694 2362
rect -2598 5150 -2316 5582
rect -2598 1930 -2316 2362
rect -2220 5150 -1938 5582
rect -2220 1930 -1938 2362
rect -1842 5150 -1560 5582
rect -1842 1930 -1560 2362
rect -1464 5150 -1182 5582
rect -1464 1930 -1182 2362
rect -1086 5150 -804 5582
rect -1086 1930 -804 2362
rect -708 5150 -426 5582
rect -708 1930 -426 2362
rect -330 5150 -48 5582
rect -330 1930 -48 2362
rect 48 5150 330 5582
rect 48 1930 330 2362
rect 426 5150 708 5582
rect 426 1930 708 2362
rect 804 5150 1086 5582
rect 804 1930 1086 2362
rect 1182 5150 1464 5582
rect 1182 1930 1464 2362
rect 1560 5150 1842 5582
rect 1560 1930 1842 2362
rect 1938 5150 2220 5582
rect 1938 1930 2220 2362
rect 2316 5150 2598 5582
rect 2316 1930 2598 2362
rect 2694 5150 2976 5582
rect 2694 1930 2976 2362
rect 3072 5150 3354 5582
rect 3072 1930 3354 2362
rect 3450 5150 3732 5582
rect 3450 1930 3732 2362
rect 3828 5150 4110 5582
rect 3828 1930 4110 2362
rect 4206 5150 4488 5582
rect 4206 1930 4488 2362
rect 4584 5150 4866 5582
rect 4584 1930 4866 2362
rect 4962 5150 5244 5582
rect 4962 1930 5244 2362
rect 5340 5150 5622 5582
rect 5340 1930 5622 2362
rect 5718 5150 6000 5582
rect 5718 1930 6000 2362
rect 6096 5150 6378 5582
rect 6096 1930 6378 2362
rect 6474 5150 6756 5582
rect 6474 1930 6756 2362
rect 6852 5150 7134 5582
rect 6852 1930 7134 2362
rect 7230 5150 7512 5582
rect 7230 1930 7512 2362
rect 7608 5150 7890 5582
rect 7608 1930 7890 2362
rect 7986 5150 8268 5582
rect 7986 1930 8268 2362
rect 8364 5150 8646 5582
rect 8364 1930 8646 2362
rect 8742 5150 9024 5582
rect 8742 1930 9024 2362
rect -9024 1394 -8742 1826
rect -9024 -1826 -8742 -1394
rect -8646 1394 -8364 1826
rect -8646 -1826 -8364 -1394
rect -8268 1394 -7986 1826
rect -8268 -1826 -7986 -1394
rect -7890 1394 -7608 1826
rect -7890 -1826 -7608 -1394
rect -7512 1394 -7230 1826
rect -7512 -1826 -7230 -1394
rect -7134 1394 -6852 1826
rect -7134 -1826 -6852 -1394
rect -6756 1394 -6474 1826
rect -6756 -1826 -6474 -1394
rect -6378 1394 -6096 1826
rect -6378 -1826 -6096 -1394
rect -6000 1394 -5718 1826
rect -6000 -1826 -5718 -1394
rect -5622 1394 -5340 1826
rect -5622 -1826 -5340 -1394
rect -5244 1394 -4962 1826
rect -5244 -1826 -4962 -1394
rect -4866 1394 -4584 1826
rect -4866 -1826 -4584 -1394
rect -4488 1394 -4206 1826
rect -4488 -1826 -4206 -1394
rect -4110 1394 -3828 1826
rect -4110 -1826 -3828 -1394
rect -3732 1394 -3450 1826
rect -3732 -1826 -3450 -1394
rect -3354 1394 -3072 1826
rect -3354 -1826 -3072 -1394
rect -2976 1394 -2694 1826
rect -2976 -1826 -2694 -1394
rect -2598 1394 -2316 1826
rect -2598 -1826 -2316 -1394
rect -2220 1394 -1938 1826
rect -2220 -1826 -1938 -1394
rect -1842 1394 -1560 1826
rect -1842 -1826 -1560 -1394
rect -1464 1394 -1182 1826
rect -1464 -1826 -1182 -1394
rect -1086 1394 -804 1826
rect -1086 -1826 -804 -1394
rect -708 1394 -426 1826
rect -708 -1826 -426 -1394
rect -330 1394 -48 1826
rect -330 -1826 -48 -1394
rect 48 1394 330 1826
rect 48 -1826 330 -1394
rect 426 1394 708 1826
rect 426 -1826 708 -1394
rect 804 1394 1086 1826
rect 804 -1826 1086 -1394
rect 1182 1394 1464 1826
rect 1182 -1826 1464 -1394
rect 1560 1394 1842 1826
rect 1560 -1826 1842 -1394
rect 1938 1394 2220 1826
rect 1938 -1826 2220 -1394
rect 2316 1394 2598 1826
rect 2316 -1826 2598 -1394
rect 2694 1394 2976 1826
rect 2694 -1826 2976 -1394
rect 3072 1394 3354 1826
rect 3072 -1826 3354 -1394
rect 3450 1394 3732 1826
rect 3450 -1826 3732 -1394
rect 3828 1394 4110 1826
rect 3828 -1826 4110 -1394
rect 4206 1394 4488 1826
rect 4206 -1826 4488 -1394
rect 4584 1394 4866 1826
rect 4584 -1826 4866 -1394
rect 4962 1394 5244 1826
rect 4962 -1826 5244 -1394
rect 5340 1394 5622 1826
rect 5340 -1826 5622 -1394
rect 5718 1394 6000 1826
rect 5718 -1826 6000 -1394
rect 6096 1394 6378 1826
rect 6096 -1826 6378 -1394
rect 6474 1394 6756 1826
rect 6474 -1826 6756 -1394
rect 6852 1394 7134 1826
rect 6852 -1826 7134 -1394
rect 7230 1394 7512 1826
rect 7230 -1826 7512 -1394
rect 7608 1394 7890 1826
rect 7608 -1826 7890 -1394
rect 7986 1394 8268 1826
rect 7986 -1826 8268 -1394
rect 8364 1394 8646 1826
rect 8364 -1826 8646 -1394
rect 8742 1394 9024 1826
rect 8742 -1826 9024 -1394
rect -9024 -2362 -8742 -1930
rect -9024 -5582 -8742 -5150
rect -8646 -2362 -8364 -1930
rect -8646 -5582 -8364 -5150
rect -8268 -2362 -7986 -1930
rect -8268 -5582 -7986 -5150
rect -7890 -2362 -7608 -1930
rect -7890 -5582 -7608 -5150
rect -7512 -2362 -7230 -1930
rect -7512 -5582 -7230 -5150
rect -7134 -2362 -6852 -1930
rect -7134 -5582 -6852 -5150
rect -6756 -2362 -6474 -1930
rect -6756 -5582 -6474 -5150
rect -6378 -2362 -6096 -1930
rect -6378 -5582 -6096 -5150
rect -6000 -2362 -5718 -1930
rect -6000 -5582 -5718 -5150
rect -5622 -2362 -5340 -1930
rect -5622 -5582 -5340 -5150
rect -5244 -2362 -4962 -1930
rect -5244 -5582 -4962 -5150
rect -4866 -2362 -4584 -1930
rect -4866 -5582 -4584 -5150
rect -4488 -2362 -4206 -1930
rect -4488 -5582 -4206 -5150
rect -4110 -2362 -3828 -1930
rect -4110 -5582 -3828 -5150
rect -3732 -2362 -3450 -1930
rect -3732 -5582 -3450 -5150
rect -3354 -2362 -3072 -1930
rect -3354 -5582 -3072 -5150
rect -2976 -2362 -2694 -1930
rect -2976 -5582 -2694 -5150
rect -2598 -2362 -2316 -1930
rect -2598 -5582 -2316 -5150
rect -2220 -2362 -1938 -1930
rect -2220 -5582 -1938 -5150
rect -1842 -2362 -1560 -1930
rect -1842 -5582 -1560 -5150
rect -1464 -2362 -1182 -1930
rect -1464 -5582 -1182 -5150
rect -1086 -2362 -804 -1930
rect -1086 -5582 -804 -5150
rect -708 -2362 -426 -1930
rect -708 -5582 -426 -5150
rect -330 -2362 -48 -1930
rect -330 -5582 -48 -5150
rect 48 -2362 330 -1930
rect 48 -5582 330 -5150
rect 426 -2362 708 -1930
rect 426 -5582 708 -5150
rect 804 -2362 1086 -1930
rect 804 -5582 1086 -5150
rect 1182 -2362 1464 -1930
rect 1182 -5582 1464 -5150
rect 1560 -2362 1842 -1930
rect 1560 -5582 1842 -5150
rect 1938 -2362 2220 -1930
rect 1938 -5582 2220 -5150
rect 2316 -2362 2598 -1930
rect 2316 -5582 2598 -5150
rect 2694 -2362 2976 -1930
rect 2694 -5582 2976 -5150
rect 3072 -2362 3354 -1930
rect 3072 -5582 3354 -5150
rect 3450 -2362 3732 -1930
rect 3450 -5582 3732 -5150
rect 3828 -2362 4110 -1930
rect 3828 -5582 4110 -5150
rect 4206 -2362 4488 -1930
rect 4206 -5582 4488 -5150
rect 4584 -2362 4866 -1930
rect 4584 -5582 4866 -5150
rect 4962 -2362 5244 -1930
rect 4962 -5582 5244 -5150
rect 5340 -2362 5622 -1930
rect 5340 -5582 5622 -5150
rect 5718 -2362 6000 -1930
rect 5718 -5582 6000 -5150
rect 6096 -2362 6378 -1930
rect 6096 -5582 6378 -5150
rect 6474 -2362 6756 -1930
rect 6474 -5582 6756 -5150
rect 6852 -2362 7134 -1930
rect 6852 -5582 7134 -5150
rect 7230 -2362 7512 -1930
rect 7230 -5582 7512 -5150
rect 7608 -2362 7890 -1930
rect 7608 -5582 7890 -5150
rect 7986 -2362 8268 -1930
rect 7986 -5582 8268 -5150
rect 8364 -2362 8646 -1930
rect 8364 -5582 8646 -5150
rect 8742 -2362 9024 -1930
rect 8742 -5582 9024 -5150
<< xpolyres >>
rect -9024 2362 -8742 5150
rect -8646 2362 -8364 5150
rect -8268 2362 -7986 5150
rect -7890 2362 -7608 5150
rect -7512 2362 -7230 5150
rect -7134 2362 -6852 5150
rect -6756 2362 -6474 5150
rect -6378 2362 -6096 5150
rect -6000 2362 -5718 5150
rect -5622 2362 -5340 5150
rect -5244 2362 -4962 5150
rect -4866 2362 -4584 5150
rect -4488 2362 -4206 5150
rect -4110 2362 -3828 5150
rect -3732 2362 -3450 5150
rect -3354 2362 -3072 5150
rect -2976 2362 -2694 5150
rect -2598 2362 -2316 5150
rect -2220 2362 -1938 5150
rect -1842 2362 -1560 5150
rect -1464 2362 -1182 5150
rect -1086 2362 -804 5150
rect -708 2362 -426 5150
rect -330 2362 -48 5150
rect 48 2362 330 5150
rect 426 2362 708 5150
rect 804 2362 1086 5150
rect 1182 2362 1464 5150
rect 1560 2362 1842 5150
rect 1938 2362 2220 5150
rect 2316 2362 2598 5150
rect 2694 2362 2976 5150
rect 3072 2362 3354 5150
rect 3450 2362 3732 5150
rect 3828 2362 4110 5150
rect 4206 2362 4488 5150
rect 4584 2362 4866 5150
rect 4962 2362 5244 5150
rect 5340 2362 5622 5150
rect 5718 2362 6000 5150
rect 6096 2362 6378 5150
rect 6474 2362 6756 5150
rect 6852 2362 7134 5150
rect 7230 2362 7512 5150
rect 7608 2362 7890 5150
rect 7986 2362 8268 5150
rect 8364 2362 8646 5150
rect 8742 2362 9024 5150
rect -9024 -1394 -8742 1394
rect -8646 -1394 -8364 1394
rect -8268 -1394 -7986 1394
rect -7890 -1394 -7608 1394
rect -7512 -1394 -7230 1394
rect -7134 -1394 -6852 1394
rect -6756 -1394 -6474 1394
rect -6378 -1394 -6096 1394
rect -6000 -1394 -5718 1394
rect -5622 -1394 -5340 1394
rect -5244 -1394 -4962 1394
rect -4866 -1394 -4584 1394
rect -4488 -1394 -4206 1394
rect -4110 -1394 -3828 1394
rect -3732 -1394 -3450 1394
rect -3354 -1394 -3072 1394
rect -2976 -1394 -2694 1394
rect -2598 -1394 -2316 1394
rect -2220 -1394 -1938 1394
rect -1842 -1394 -1560 1394
rect -1464 -1394 -1182 1394
rect -1086 -1394 -804 1394
rect -708 -1394 -426 1394
rect -330 -1394 -48 1394
rect 48 -1394 330 1394
rect 426 -1394 708 1394
rect 804 -1394 1086 1394
rect 1182 -1394 1464 1394
rect 1560 -1394 1842 1394
rect 1938 -1394 2220 1394
rect 2316 -1394 2598 1394
rect 2694 -1394 2976 1394
rect 3072 -1394 3354 1394
rect 3450 -1394 3732 1394
rect 3828 -1394 4110 1394
rect 4206 -1394 4488 1394
rect 4584 -1394 4866 1394
rect 4962 -1394 5244 1394
rect 5340 -1394 5622 1394
rect 5718 -1394 6000 1394
rect 6096 -1394 6378 1394
rect 6474 -1394 6756 1394
rect 6852 -1394 7134 1394
rect 7230 -1394 7512 1394
rect 7608 -1394 7890 1394
rect 7986 -1394 8268 1394
rect 8364 -1394 8646 1394
rect 8742 -1394 9024 1394
rect -9024 -5150 -8742 -2362
rect -8646 -5150 -8364 -2362
rect -8268 -5150 -7986 -2362
rect -7890 -5150 -7608 -2362
rect -7512 -5150 -7230 -2362
rect -7134 -5150 -6852 -2362
rect -6756 -5150 -6474 -2362
rect -6378 -5150 -6096 -2362
rect -6000 -5150 -5718 -2362
rect -5622 -5150 -5340 -2362
rect -5244 -5150 -4962 -2362
rect -4866 -5150 -4584 -2362
rect -4488 -5150 -4206 -2362
rect -4110 -5150 -3828 -2362
rect -3732 -5150 -3450 -2362
rect -3354 -5150 -3072 -2362
rect -2976 -5150 -2694 -2362
rect -2598 -5150 -2316 -2362
rect -2220 -5150 -1938 -2362
rect -1842 -5150 -1560 -2362
rect -1464 -5150 -1182 -2362
rect -1086 -5150 -804 -2362
rect -708 -5150 -426 -2362
rect -330 -5150 -48 -2362
rect 48 -5150 330 -2362
rect 426 -5150 708 -2362
rect 804 -5150 1086 -2362
rect 1182 -5150 1464 -2362
rect 1560 -5150 1842 -2362
rect 1938 -5150 2220 -2362
rect 2316 -5150 2598 -2362
rect 2694 -5150 2976 -2362
rect 3072 -5150 3354 -2362
rect 3450 -5150 3732 -2362
rect 3828 -5150 4110 -2362
rect 4206 -5150 4488 -2362
rect 4584 -5150 4866 -2362
rect 4962 -5150 5244 -2362
rect 5340 -5150 5622 -2362
rect 5718 -5150 6000 -2362
rect 6096 -5150 6378 -2362
rect 6474 -5150 6756 -2362
rect 6852 -5150 7134 -2362
rect 7230 -5150 7512 -2362
rect 7608 -5150 7890 -2362
rect 7986 -5150 8268 -2362
rect 8364 -5150 8646 -2362
rect 8742 -5150 9024 -2362
<< viali >>
rect -9008 5167 -8758 5564
rect -8630 5167 -8380 5564
rect -8252 5167 -8002 5564
rect -7874 5167 -7624 5564
rect -7496 5167 -7246 5564
rect -7118 5167 -6868 5564
rect -6740 5167 -6490 5564
rect -6362 5167 -6112 5564
rect -5984 5167 -5734 5564
rect -5606 5167 -5356 5564
rect -5228 5167 -4978 5564
rect -4850 5167 -4600 5564
rect -4472 5167 -4222 5564
rect -4094 5167 -3844 5564
rect -3716 5167 -3466 5564
rect -3338 5167 -3088 5564
rect -2960 5167 -2710 5564
rect -2582 5167 -2332 5564
rect -2204 5167 -1954 5564
rect -1826 5167 -1576 5564
rect -1448 5167 -1198 5564
rect -1070 5167 -820 5564
rect -692 5167 -442 5564
rect -314 5167 -64 5564
rect 64 5167 314 5564
rect 442 5167 692 5564
rect 820 5167 1070 5564
rect 1198 5167 1448 5564
rect 1576 5167 1826 5564
rect 1954 5167 2204 5564
rect 2332 5167 2582 5564
rect 2710 5167 2960 5564
rect 3088 5167 3338 5564
rect 3466 5167 3716 5564
rect 3844 5167 4094 5564
rect 4222 5167 4472 5564
rect 4600 5167 4850 5564
rect 4978 5167 5228 5564
rect 5356 5167 5606 5564
rect 5734 5167 5984 5564
rect 6112 5167 6362 5564
rect 6490 5167 6740 5564
rect 6868 5167 7118 5564
rect 7246 5167 7496 5564
rect 7624 5167 7874 5564
rect 8002 5167 8252 5564
rect 8380 5167 8630 5564
rect 8758 5167 9008 5564
rect -9008 1948 -8758 2345
rect -8630 1948 -8380 2345
rect -8252 1948 -8002 2345
rect -7874 1948 -7624 2345
rect -7496 1948 -7246 2345
rect -7118 1948 -6868 2345
rect -6740 1948 -6490 2345
rect -6362 1948 -6112 2345
rect -5984 1948 -5734 2345
rect -5606 1948 -5356 2345
rect -5228 1948 -4978 2345
rect -4850 1948 -4600 2345
rect -4472 1948 -4222 2345
rect -4094 1948 -3844 2345
rect -3716 1948 -3466 2345
rect -3338 1948 -3088 2345
rect -2960 1948 -2710 2345
rect -2582 1948 -2332 2345
rect -2204 1948 -1954 2345
rect -1826 1948 -1576 2345
rect -1448 1948 -1198 2345
rect -1070 1948 -820 2345
rect -692 1948 -442 2345
rect -314 1948 -64 2345
rect 64 1948 314 2345
rect 442 1948 692 2345
rect 820 1948 1070 2345
rect 1198 1948 1448 2345
rect 1576 1948 1826 2345
rect 1954 1948 2204 2345
rect 2332 1948 2582 2345
rect 2710 1948 2960 2345
rect 3088 1948 3338 2345
rect 3466 1948 3716 2345
rect 3844 1948 4094 2345
rect 4222 1948 4472 2345
rect 4600 1948 4850 2345
rect 4978 1948 5228 2345
rect 5356 1948 5606 2345
rect 5734 1948 5984 2345
rect 6112 1948 6362 2345
rect 6490 1948 6740 2345
rect 6868 1948 7118 2345
rect 7246 1948 7496 2345
rect 7624 1948 7874 2345
rect 8002 1948 8252 2345
rect 8380 1948 8630 2345
rect 8758 1948 9008 2345
rect -9008 1411 -8758 1808
rect -8630 1411 -8380 1808
rect -8252 1411 -8002 1808
rect -7874 1411 -7624 1808
rect -7496 1411 -7246 1808
rect -7118 1411 -6868 1808
rect -6740 1411 -6490 1808
rect -6362 1411 -6112 1808
rect -5984 1411 -5734 1808
rect -5606 1411 -5356 1808
rect -5228 1411 -4978 1808
rect -4850 1411 -4600 1808
rect -4472 1411 -4222 1808
rect -4094 1411 -3844 1808
rect -3716 1411 -3466 1808
rect -3338 1411 -3088 1808
rect -2960 1411 -2710 1808
rect -2582 1411 -2332 1808
rect -2204 1411 -1954 1808
rect -1826 1411 -1576 1808
rect -1448 1411 -1198 1808
rect -1070 1411 -820 1808
rect -692 1411 -442 1808
rect -314 1411 -64 1808
rect 64 1411 314 1808
rect 442 1411 692 1808
rect 820 1411 1070 1808
rect 1198 1411 1448 1808
rect 1576 1411 1826 1808
rect 1954 1411 2204 1808
rect 2332 1411 2582 1808
rect 2710 1411 2960 1808
rect 3088 1411 3338 1808
rect 3466 1411 3716 1808
rect 3844 1411 4094 1808
rect 4222 1411 4472 1808
rect 4600 1411 4850 1808
rect 4978 1411 5228 1808
rect 5356 1411 5606 1808
rect 5734 1411 5984 1808
rect 6112 1411 6362 1808
rect 6490 1411 6740 1808
rect 6868 1411 7118 1808
rect 7246 1411 7496 1808
rect 7624 1411 7874 1808
rect 8002 1411 8252 1808
rect 8380 1411 8630 1808
rect 8758 1411 9008 1808
rect -9008 -1808 -8758 -1411
rect -8630 -1808 -8380 -1411
rect -8252 -1808 -8002 -1411
rect -7874 -1808 -7624 -1411
rect -7496 -1808 -7246 -1411
rect -7118 -1808 -6868 -1411
rect -6740 -1808 -6490 -1411
rect -6362 -1808 -6112 -1411
rect -5984 -1808 -5734 -1411
rect -5606 -1808 -5356 -1411
rect -5228 -1808 -4978 -1411
rect -4850 -1808 -4600 -1411
rect -4472 -1808 -4222 -1411
rect -4094 -1808 -3844 -1411
rect -3716 -1808 -3466 -1411
rect -3338 -1808 -3088 -1411
rect -2960 -1808 -2710 -1411
rect -2582 -1808 -2332 -1411
rect -2204 -1808 -1954 -1411
rect -1826 -1808 -1576 -1411
rect -1448 -1808 -1198 -1411
rect -1070 -1808 -820 -1411
rect -692 -1808 -442 -1411
rect -314 -1808 -64 -1411
rect 64 -1808 314 -1411
rect 442 -1808 692 -1411
rect 820 -1808 1070 -1411
rect 1198 -1808 1448 -1411
rect 1576 -1808 1826 -1411
rect 1954 -1808 2204 -1411
rect 2332 -1808 2582 -1411
rect 2710 -1808 2960 -1411
rect 3088 -1808 3338 -1411
rect 3466 -1808 3716 -1411
rect 3844 -1808 4094 -1411
rect 4222 -1808 4472 -1411
rect 4600 -1808 4850 -1411
rect 4978 -1808 5228 -1411
rect 5356 -1808 5606 -1411
rect 5734 -1808 5984 -1411
rect 6112 -1808 6362 -1411
rect 6490 -1808 6740 -1411
rect 6868 -1808 7118 -1411
rect 7246 -1808 7496 -1411
rect 7624 -1808 7874 -1411
rect 8002 -1808 8252 -1411
rect 8380 -1808 8630 -1411
rect 8758 -1808 9008 -1411
rect -9008 -2345 -8758 -1948
rect -8630 -2345 -8380 -1948
rect -8252 -2345 -8002 -1948
rect -7874 -2345 -7624 -1948
rect -7496 -2345 -7246 -1948
rect -7118 -2345 -6868 -1948
rect -6740 -2345 -6490 -1948
rect -6362 -2345 -6112 -1948
rect -5984 -2345 -5734 -1948
rect -5606 -2345 -5356 -1948
rect -5228 -2345 -4978 -1948
rect -4850 -2345 -4600 -1948
rect -4472 -2345 -4222 -1948
rect -4094 -2345 -3844 -1948
rect -3716 -2345 -3466 -1948
rect -3338 -2345 -3088 -1948
rect -2960 -2345 -2710 -1948
rect -2582 -2345 -2332 -1948
rect -2204 -2345 -1954 -1948
rect -1826 -2345 -1576 -1948
rect -1448 -2345 -1198 -1948
rect -1070 -2345 -820 -1948
rect -692 -2345 -442 -1948
rect -314 -2345 -64 -1948
rect 64 -2345 314 -1948
rect 442 -2345 692 -1948
rect 820 -2345 1070 -1948
rect 1198 -2345 1448 -1948
rect 1576 -2345 1826 -1948
rect 1954 -2345 2204 -1948
rect 2332 -2345 2582 -1948
rect 2710 -2345 2960 -1948
rect 3088 -2345 3338 -1948
rect 3466 -2345 3716 -1948
rect 3844 -2345 4094 -1948
rect 4222 -2345 4472 -1948
rect 4600 -2345 4850 -1948
rect 4978 -2345 5228 -1948
rect 5356 -2345 5606 -1948
rect 5734 -2345 5984 -1948
rect 6112 -2345 6362 -1948
rect 6490 -2345 6740 -1948
rect 6868 -2345 7118 -1948
rect 7246 -2345 7496 -1948
rect 7624 -2345 7874 -1948
rect 8002 -2345 8252 -1948
rect 8380 -2345 8630 -1948
rect 8758 -2345 9008 -1948
rect -9008 -5564 -8758 -5167
rect -8630 -5564 -8380 -5167
rect -8252 -5564 -8002 -5167
rect -7874 -5564 -7624 -5167
rect -7496 -5564 -7246 -5167
rect -7118 -5564 -6868 -5167
rect -6740 -5564 -6490 -5167
rect -6362 -5564 -6112 -5167
rect -5984 -5564 -5734 -5167
rect -5606 -5564 -5356 -5167
rect -5228 -5564 -4978 -5167
rect -4850 -5564 -4600 -5167
rect -4472 -5564 -4222 -5167
rect -4094 -5564 -3844 -5167
rect -3716 -5564 -3466 -5167
rect -3338 -5564 -3088 -5167
rect -2960 -5564 -2710 -5167
rect -2582 -5564 -2332 -5167
rect -2204 -5564 -1954 -5167
rect -1826 -5564 -1576 -5167
rect -1448 -5564 -1198 -5167
rect -1070 -5564 -820 -5167
rect -692 -5564 -442 -5167
rect -314 -5564 -64 -5167
rect 64 -5564 314 -5167
rect 442 -5564 692 -5167
rect 820 -5564 1070 -5167
rect 1198 -5564 1448 -5167
rect 1576 -5564 1826 -5167
rect 1954 -5564 2204 -5167
rect 2332 -5564 2582 -5167
rect 2710 -5564 2960 -5167
rect 3088 -5564 3338 -5167
rect 3466 -5564 3716 -5167
rect 3844 -5564 4094 -5167
rect 4222 -5564 4472 -5167
rect 4600 -5564 4850 -5167
rect 4978 -5564 5228 -5167
rect 5356 -5564 5606 -5167
rect 5734 -5564 5984 -5167
rect 6112 -5564 6362 -5167
rect 6490 -5564 6740 -5167
rect 6868 -5564 7118 -5167
rect 7246 -5564 7496 -5167
rect 7624 -5564 7874 -5167
rect 8002 -5564 8252 -5167
rect 8380 -5564 8630 -5167
rect 8758 -5564 9008 -5167
<< metal1 >>
rect -9014 5564 -8752 5576
rect -9014 5167 -9008 5564
rect -8758 5167 -8752 5564
rect -9014 5155 -8752 5167
rect -8636 5564 -8374 5576
rect -8636 5167 -8630 5564
rect -8380 5167 -8374 5564
rect -8636 5155 -8374 5167
rect -8258 5564 -7996 5576
rect -8258 5167 -8252 5564
rect -8002 5167 -7996 5564
rect -8258 5155 -7996 5167
rect -7880 5564 -7618 5576
rect -7880 5167 -7874 5564
rect -7624 5167 -7618 5564
rect -7880 5155 -7618 5167
rect -7502 5564 -7240 5576
rect -7502 5167 -7496 5564
rect -7246 5167 -7240 5564
rect -7502 5155 -7240 5167
rect -7124 5564 -6862 5576
rect -7124 5167 -7118 5564
rect -6868 5167 -6862 5564
rect -7124 5155 -6862 5167
rect -6746 5564 -6484 5576
rect -6746 5167 -6740 5564
rect -6490 5167 -6484 5564
rect -6746 5155 -6484 5167
rect -6368 5564 -6106 5576
rect -6368 5167 -6362 5564
rect -6112 5167 -6106 5564
rect -6368 5155 -6106 5167
rect -5990 5564 -5728 5576
rect -5990 5167 -5984 5564
rect -5734 5167 -5728 5564
rect -5990 5155 -5728 5167
rect -5612 5564 -5350 5576
rect -5612 5167 -5606 5564
rect -5356 5167 -5350 5564
rect -5612 5155 -5350 5167
rect -5234 5564 -4972 5576
rect -5234 5167 -5228 5564
rect -4978 5167 -4972 5564
rect -5234 5155 -4972 5167
rect -4856 5564 -4594 5576
rect -4856 5167 -4850 5564
rect -4600 5167 -4594 5564
rect -4856 5155 -4594 5167
rect -4478 5564 -4216 5576
rect -4478 5167 -4472 5564
rect -4222 5167 -4216 5564
rect -4478 5155 -4216 5167
rect -4100 5564 -3838 5576
rect -4100 5167 -4094 5564
rect -3844 5167 -3838 5564
rect -4100 5155 -3838 5167
rect -3722 5564 -3460 5576
rect -3722 5167 -3716 5564
rect -3466 5167 -3460 5564
rect -3722 5155 -3460 5167
rect -3344 5564 -3082 5576
rect -3344 5167 -3338 5564
rect -3088 5167 -3082 5564
rect -3344 5155 -3082 5167
rect -2966 5564 -2704 5576
rect -2966 5167 -2960 5564
rect -2710 5167 -2704 5564
rect -2966 5155 -2704 5167
rect -2588 5564 -2326 5576
rect -2588 5167 -2582 5564
rect -2332 5167 -2326 5564
rect -2588 5155 -2326 5167
rect -2210 5564 -1948 5576
rect -2210 5167 -2204 5564
rect -1954 5167 -1948 5564
rect -2210 5155 -1948 5167
rect -1832 5564 -1570 5576
rect -1832 5167 -1826 5564
rect -1576 5167 -1570 5564
rect -1832 5155 -1570 5167
rect -1454 5564 -1192 5576
rect -1454 5167 -1448 5564
rect -1198 5167 -1192 5564
rect -1454 5155 -1192 5167
rect -1076 5564 -814 5576
rect -1076 5167 -1070 5564
rect -820 5167 -814 5564
rect -1076 5155 -814 5167
rect -698 5564 -436 5576
rect -698 5167 -692 5564
rect -442 5167 -436 5564
rect -698 5155 -436 5167
rect -320 5564 -58 5576
rect -320 5167 -314 5564
rect -64 5167 -58 5564
rect -320 5155 -58 5167
rect 58 5564 320 5576
rect 58 5167 64 5564
rect 314 5167 320 5564
rect 58 5155 320 5167
rect 436 5564 698 5576
rect 436 5167 442 5564
rect 692 5167 698 5564
rect 436 5155 698 5167
rect 814 5564 1076 5576
rect 814 5167 820 5564
rect 1070 5167 1076 5564
rect 814 5155 1076 5167
rect 1192 5564 1454 5576
rect 1192 5167 1198 5564
rect 1448 5167 1454 5564
rect 1192 5155 1454 5167
rect 1570 5564 1832 5576
rect 1570 5167 1576 5564
rect 1826 5167 1832 5564
rect 1570 5155 1832 5167
rect 1948 5564 2210 5576
rect 1948 5167 1954 5564
rect 2204 5167 2210 5564
rect 1948 5155 2210 5167
rect 2326 5564 2588 5576
rect 2326 5167 2332 5564
rect 2582 5167 2588 5564
rect 2326 5155 2588 5167
rect 2704 5564 2966 5576
rect 2704 5167 2710 5564
rect 2960 5167 2966 5564
rect 2704 5155 2966 5167
rect 3082 5564 3344 5576
rect 3082 5167 3088 5564
rect 3338 5167 3344 5564
rect 3082 5155 3344 5167
rect 3460 5564 3722 5576
rect 3460 5167 3466 5564
rect 3716 5167 3722 5564
rect 3460 5155 3722 5167
rect 3838 5564 4100 5576
rect 3838 5167 3844 5564
rect 4094 5167 4100 5564
rect 3838 5155 4100 5167
rect 4216 5564 4478 5576
rect 4216 5167 4222 5564
rect 4472 5167 4478 5564
rect 4216 5155 4478 5167
rect 4594 5564 4856 5576
rect 4594 5167 4600 5564
rect 4850 5167 4856 5564
rect 4594 5155 4856 5167
rect 4972 5564 5234 5576
rect 4972 5167 4978 5564
rect 5228 5167 5234 5564
rect 4972 5155 5234 5167
rect 5350 5564 5612 5576
rect 5350 5167 5356 5564
rect 5606 5167 5612 5564
rect 5350 5155 5612 5167
rect 5728 5564 5990 5576
rect 5728 5167 5734 5564
rect 5984 5167 5990 5564
rect 5728 5155 5990 5167
rect 6106 5564 6368 5576
rect 6106 5167 6112 5564
rect 6362 5167 6368 5564
rect 6106 5155 6368 5167
rect 6484 5564 6746 5576
rect 6484 5167 6490 5564
rect 6740 5167 6746 5564
rect 6484 5155 6746 5167
rect 6862 5564 7124 5576
rect 6862 5167 6868 5564
rect 7118 5167 7124 5564
rect 6862 5155 7124 5167
rect 7240 5564 7502 5576
rect 7240 5167 7246 5564
rect 7496 5167 7502 5564
rect 7240 5155 7502 5167
rect 7618 5564 7880 5576
rect 7618 5167 7624 5564
rect 7874 5167 7880 5564
rect 7618 5155 7880 5167
rect 7996 5564 8258 5576
rect 7996 5167 8002 5564
rect 8252 5167 8258 5564
rect 7996 5155 8258 5167
rect 8374 5564 8636 5576
rect 8374 5167 8380 5564
rect 8630 5167 8636 5564
rect 8374 5155 8636 5167
rect 8752 5564 9014 5576
rect 8752 5167 8758 5564
rect 9008 5167 9014 5564
rect 8752 5155 9014 5167
rect -9014 2345 -8752 2357
rect -9014 1948 -9008 2345
rect -8758 1948 -8752 2345
rect -9014 1936 -8752 1948
rect -8636 2345 -8374 2357
rect -8636 1948 -8630 2345
rect -8380 1948 -8374 2345
rect -8636 1936 -8374 1948
rect -8258 2345 -7996 2357
rect -8258 1948 -8252 2345
rect -8002 1948 -7996 2345
rect -8258 1936 -7996 1948
rect -7880 2345 -7618 2357
rect -7880 1948 -7874 2345
rect -7624 1948 -7618 2345
rect -7880 1936 -7618 1948
rect -7502 2345 -7240 2357
rect -7502 1948 -7496 2345
rect -7246 1948 -7240 2345
rect -7502 1936 -7240 1948
rect -7124 2345 -6862 2357
rect -7124 1948 -7118 2345
rect -6868 1948 -6862 2345
rect -7124 1936 -6862 1948
rect -6746 2345 -6484 2357
rect -6746 1948 -6740 2345
rect -6490 1948 -6484 2345
rect -6746 1936 -6484 1948
rect -6368 2345 -6106 2357
rect -6368 1948 -6362 2345
rect -6112 1948 -6106 2345
rect -6368 1936 -6106 1948
rect -5990 2345 -5728 2357
rect -5990 1948 -5984 2345
rect -5734 1948 -5728 2345
rect -5990 1936 -5728 1948
rect -5612 2345 -5350 2357
rect -5612 1948 -5606 2345
rect -5356 1948 -5350 2345
rect -5612 1936 -5350 1948
rect -5234 2345 -4972 2357
rect -5234 1948 -5228 2345
rect -4978 1948 -4972 2345
rect -5234 1936 -4972 1948
rect -4856 2345 -4594 2357
rect -4856 1948 -4850 2345
rect -4600 1948 -4594 2345
rect -4856 1936 -4594 1948
rect -4478 2345 -4216 2357
rect -4478 1948 -4472 2345
rect -4222 1948 -4216 2345
rect -4478 1936 -4216 1948
rect -4100 2345 -3838 2357
rect -4100 1948 -4094 2345
rect -3844 1948 -3838 2345
rect -4100 1936 -3838 1948
rect -3722 2345 -3460 2357
rect -3722 1948 -3716 2345
rect -3466 1948 -3460 2345
rect -3722 1936 -3460 1948
rect -3344 2345 -3082 2357
rect -3344 1948 -3338 2345
rect -3088 1948 -3082 2345
rect -3344 1936 -3082 1948
rect -2966 2345 -2704 2357
rect -2966 1948 -2960 2345
rect -2710 1948 -2704 2345
rect -2966 1936 -2704 1948
rect -2588 2345 -2326 2357
rect -2588 1948 -2582 2345
rect -2332 1948 -2326 2345
rect -2588 1936 -2326 1948
rect -2210 2345 -1948 2357
rect -2210 1948 -2204 2345
rect -1954 1948 -1948 2345
rect -2210 1936 -1948 1948
rect -1832 2345 -1570 2357
rect -1832 1948 -1826 2345
rect -1576 1948 -1570 2345
rect -1832 1936 -1570 1948
rect -1454 2345 -1192 2357
rect -1454 1948 -1448 2345
rect -1198 1948 -1192 2345
rect -1454 1936 -1192 1948
rect -1076 2345 -814 2357
rect -1076 1948 -1070 2345
rect -820 1948 -814 2345
rect -1076 1936 -814 1948
rect -698 2345 -436 2357
rect -698 1948 -692 2345
rect -442 1948 -436 2345
rect -698 1936 -436 1948
rect -320 2345 -58 2357
rect -320 1948 -314 2345
rect -64 1948 -58 2345
rect -320 1936 -58 1948
rect 58 2345 320 2357
rect 58 1948 64 2345
rect 314 1948 320 2345
rect 58 1936 320 1948
rect 436 2345 698 2357
rect 436 1948 442 2345
rect 692 1948 698 2345
rect 436 1936 698 1948
rect 814 2345 1076 2357
rect 814 1948 820 2345
rect 1070 1948 1076 2345
rect 814 1936 1076 1948
rect 1192 2345 1454 2357
rect 1192 1948 1198 2345
rect 1448 1948 1454 2345
rect 1192 1936 1454 1948
rect 1570 2345 1832 2357
rect 1570 1948 1576 2345
rect 1826 1948 1832 2345
rect 1570 1936 1832 1948
rect 1948 2345 2210 2357
rect 1948 1948 1954 2345
rect 2204 1948 2210 2345
rect 1948 1936 2210 1948
rect 2326 2345 2588 2357
rect 2326 1948 2332 2345
rect 2582 1948 2588 2345
rect 2326 1936 2588 1948
rect 2704 2345 2966 2357
rect 2704 1948 2710 2345
rect 2960 1948 2966 2345
rect 2704 1936 2966 1948
rect 3082 2345 3344 2357
rect 3082 1948 3088 2345
rect 3338 1948 3344 2345
rect 3082 1936 3344 1948
rect 3460 2345 3722 2357
rect 3460 1948 3466 2345
rect 3716 1948 3722 2345
rect 3460 1936 3722 1948
rect 3838 2345 4100 2357
rect 3838 1948 3844 2345
rect 4094 1948 4100 2345
rect 3838 1936 4100 1948
rect 4216 2345 4478 2357
rect 4216 1948 4222 2345
rect 4472 1948 4478 2345
rect 4216 1936 4478 1948
rect 4594 2345 4856 2357
rect 4594 1948 4600 2345
rect 4850 1948 4856 2345
rect 4594 1936 4856 1948
rect 4972 2345 5234 2357
rect 4972 1948 4978 2345
rect 5228 1948 5234 2345
rect 4972 1936 5234 1948
rect 5350 2345 5612 2357
rect 5350 1948 5356 2345
rect 5606 1948 5612 2345
rect 5350 1936 5612 1948
rect 5728 2345 5990 2357
rect 5728 1948 5734 2345
rect 5984 1948 5990 2345
rect 5728 1936 5990 1948
rect 6106 2345 6368 2357
rect 6106 1948 6112 2345
rect 6362 1948 6368 2345
rect 6106 1936 6368 1948
rect 6484 2345 6746 2357
rect 6484 1948 6490 2345
rect 6740 1948 6746 2345
rect 6484 1936 6746 1948
rect 6862 2345 7124 2357
rect 6862 1948 6868 2345
rect 7118 1948 7124 2345
rect 6862 1936 7124 1948
rect 7240 2345 7502 2357
rect 7240 1948 7246 2345
rect 7496 1948 7502 2345
rect 7240 1936 7502 1948
rect 7618 2345 7880 2357
rect 7618 1948 7624 2345
rect 7874 1948 7880 2345
rect 7618 1936 7880 1948
rect 7996 2345 8258 2357
rect 7996 1948 8002 2345
rect 8252 1948 8258 2345
rect 7996 1936 8258 1948
rect 8374 2345 8636 2357
rect 8374 1948 8380 2345
rect 8630 1948 8636 2345
rect 8374 1936 8636 1948
rect 8752 2345 9014 2357
rect 8752 1948 8758 2345
rect 9008 1948 9014 2345
rect 8752 1936 9014 1948
rect -9014 1808 -8752 1820
rect -9014 1411 -9008 1808
rect -8758 1411 -8752 1808
rect -9014 1399 -8752 1411
rect -8636 1808 -8374 1820
rect -8636 1411 -8630 1808
rect -8380 1411 -8374 1808
rect -8636 1399 -8374 1411
rect -8258 1808 -7996 1820
rect -8258 1411 -8252 1808
rect -8002 1411 -7996 1808
rect -8258 1399 -7996 1411
rect -7880 1808 -7618 1820
rect -7880 1411 -7874 1808
rect -7624 1411 -7618 1808
rect -7880 1399 -7618 1411
rect -7502 1808 -7240 1820
rect -7502 1411 -7496 1808
rect -7246 1411 -7240 1808
rect -7502 1399 -7240 1411
rect -7124 1808 -6862 1820
rect -7124 1411 -7118 1808
rect -6868 1411 -6862 1808
rect -7124 1399 -6862 1411
rect -6746 1808 -6484 1820
rect -6746 1411 -6740 1808
rect -6490 1411 -6484 1808
rect -6746 1399 -6484 1411
rect -6368 1808 -6106 1820
rect -6368 1411 -6362 1808
rect -6112 1411 -6106 1808
rect -6368 1399 -6106 1411
rect -5990 1808 -5728 1820
rect -5990 1411 -5984 1808
rect -5734 1411 -5728 1808
rect -5990 1399 -5728 1411
rect -5612 1808 -5350 1820
rect -5612 1411 -5606 1808
rect -5356 1411 -5350 1808
rect -5612 1399 -5350 1411
rect -5234 1808 -4972 1820
rect -5234 1411 -5228 1808
rect -4978 1411 -4972 1808
rect -5234 1399 -4972 1411
rect -4856 1808 -4594 1820
rect -4856 1411 -4850 1808
rect -4600 1411 -4594 1808
rect -4856 1399 -4594 1411
rect -4478 1808 -4216 1820
rect -4478 1411 -4472 1808
rect -4222 1411 -4216 1808
rect -4478 1399 -4216 1411
rect -4100 1808 -3838 1820
rect -4100 1411 -4094 1808
rect -3844 1411 -3838 1808
rect -4100 1399 -3838 1411
rect -3722 1808 -3460 1820
rect -3722 1411 -3716 1808
rect -3466 1411 -3460 1808
rect -3722 1399 -3460 1411
rect -3344 1808 -3082 1820
rect -3344 1411 -3338 1808
rect -3088 1411 -3082 1808
rect -3344 1399 -3082 1411
rect -2966 1808 -2704 1820
rect -2966 1411 -2960 1808
rect -2710 1411 -2704 1808
rect -2966 1399 -2704 1411
rect -2588 1808 -2326 1820
rect -2588 1411 -2582 1808
rect -2332 1411 -2326 1808
rect -2588 1399 -2326 1411
rect -2210 1808 -1948 1820
rect -2210 1411 -2204 1808
rect -1954 1411 -1948 1808
rect -2210 1399 -1948 1411
rect -1832 1808 -1570 1820
rect -1832 1411 -1826 1808
rect -1576 1411 -1570 1808
rect -1832 1399 -1570 1411
rect -1454 1808 -1192 1820
rect -1454 1411 -1448 1808
rect -1198 1411 -1192 1808
rect -1454 1399 -1192 1411
rect -1076 1808 -814 1820
rect -1076 1411 -1070 1808
rect -820 1411 -814 1808
rect -1076 1399 -814 1411
rect -698 1808 -436 1820
rect -698 1411 -692 1808
rect -442 1411 -436 1808
rect -698 1399 -436 1411
rect -320 1808 -58 1820
rect -320 1411 -314 1808
rect -64 1411 -58 1808
rect -320 1399 -58 1411
rect 58 1808 320 1820
rect 58 1411 64 1808
rect 314 1411 320 1808
rect 58 1399 320 1411
rect 436 1808 698 1820
rect 436 1411 442 1808
rect 692 1411 698 1808
rect 436 1399 698 1411
rect 814 1808 1076 1820
rect 814 1411 820 1808
rect 1070 1411 1076 1808
rect 814 1399 1076 1411
rect 1192 1808 1454 1820
rect 1192 1411 1198 1808
rect 1448 1411 1454 1808
rect 1192 1399 1454 1411
rect 1570 1808 1832 1820
rect 1570 1411 1576 1808
rect 1826 1411 1832 1808
rect 1570 1399 1832 1411
rect 1948 1808 2210 1820
rect 1948 1411 1954 1808
rect 2204 1411 2210 1808
rect 1948 1399 2210 1411
rect 2326 1808 2588 1820
rect 2326 1411 2332 1808
rect 2582 1411 2588 1808
rect 2326 1399 2588 1411
rect 2704 1808 2966 1820
rect 2704 1411 2710 1808
rect 2960 1411 2966 1808
rect 2704 1399 2966 1411
rect 3082 1808 3344 1820
rect 3082 1411 3088 1808
rect 3338 1411 3344 1808
rect 3082 1399 3344 1411
rect 3460 1808 3722 1820
rect 3460 1411 3466 1808
rect 3716 1411 3722 1808
rect 3460 1399 3722 1411
rect 3838 1808 4100 1820
rect 3838 1411 3844 1808
rect 4094 1411 4100 1808
rect 3838 1399 4100 1411
rect 4216 1808 4478 1820
rect 4216 1411 4222 1808
rect 4472 1411 4478 1808
rect 4216 1399 4478 1411
rect 4594 1808 4856 1820
rect 4594 1411 4600 1808
rect 4850 1411 4856 1808
rect 4594 1399 4856 1411
rect 4972 1808 5234 1820
rect 4972 1411 4978 1808
rect 5228 1411 5234 1808
rect 4972 1399 5234 1411
rect 5350 1808 5612 1820
rect 5350 1411 5356 1808
rect 5606 1411 5612 1808
rect 5350 1399 5612 1411
rect 5728 1808 5990 1820
rect 5728 1411 5734 1808
rect 5984 1411 5990 1808
rect 5728 1399 5990 1411
rect 6106 1808 6368 1820
rect 6106 1411 6112 1808
rect 6362 1411 6368 1808
rect 6106 1399 6368 1411
rect 6484 1808 6746 1820
rect 6484 1411 6490 1808
rect 6740 1411 6746 1808
rect 6484 1399 6746 1411
rect 6862 1808 7124 1820
rect 6862 1411 6868 1808
rect 7118 1411 7124 1808
rect 6862 1399 7124 1411
rect 7240 1808 7502 1820
rect 7240 1411 7246 1808
rect 7496 1411 7502 1808
rect 7240 1399 7502 1411
rect 7618 1808 7880 1820
rect 7618 1411 7624 1808
rect 7874 1411 7880 1808
rect 7618 1399 7880 1411
rect 7996 1808 8258 1820
rect 7996 1411 8002 1808
rect 8252 1411 8258 1808
rect 7996 1399 8258 1411
rect 8374 1808 8636 1820
rect 8374 1411 8380 1808
rect 8630 1411 8636 1808
rect 8374 1399 8636 1411
rect 8752 1808 9014 1820
rect 8752 1411 8758 1808
rect 9008 1411 9014 1808
rect 8752 1399 9014 1411
rect -9014 -1411 -8752 -1399
rect -9014 -1808 -9008 -1411
rect -8758 -1808 -8752 -1411
rect -9014 -1820 -8752 -1808
rect -8636 -1411 -8374 -1399
rect -8636 -1808 -8630 -1411
rect -8380 -1808 -8374 -1411
rect -8636 -1820 -8374 -1808
rect -8258 -1411 -7996 -1399
rect -8258 -1808 -8252 -1411
rect -8002 -1808 -7996 -1411
rect -8258 -1820 -7996 -1808
rect -7880 -1411 -7618 -1399
rect -7880 -1808 -7874 -1411
rect -7624 -1808 -7618 -1411
rect -7880 -1820 -7618 -1808
rect -7502 -1411 -7240 -1399
rect -7502 -1808 -7496 -1411
rect -7246 -1808 -7240 -1411
rect -7502 -1820 -7240 -1808
rect -7124 -1411 -6862 -1399
rect -7124 -1808 -7118 -1411
rect -6868 -1808 -6862 -1411
rect -7124 -1820 -6862 -1808
rect -6746 -1411 -6484 -1399
rect -6746 -1808 -6740 -1411
rect -6490 -1808 -6484 -1411
rect -6746 -1820 -6484 -1808
rect -6368 -1411 -6106 -1399
rect -6368 -1808 -6362 -1411
rect -6112 -1808 -6106 -1411
rect -6368 -1820 -6106 -1808
rect -5990 -1411 -5728 -1399
rect -5990 -1808 -5984 -1411
rect -5734 -1808 -5728 -1411
rect -5990 -1820 -5728 -1808
rect -5612 -1411 -5350 -1399
rect -5612 -1808 -5606 -1411
rect -5356 -1808 -5350 -1411
rect -5612 -1820 -5350 -1808
rect -5234 -1411 -4972 -1399
rect -5234 -1808 -5228 -1411
rect -4978 -1808 -4972 -1411
rect -5234 -1820 -4972 -1808
rect -4856 -1411 -4594 -1399
rect -4856 -1808 -4850 -1411
rect -4600 -1808 -4594 -1411
rect -4856 -1820 -4594 -1808
rect -4478 -1411 -4216 -1399
rect -4478 -1808 -4472 -1411
rect -4222 -1808 -4216 -1411
rect -4478 -1820 -4216 -1808
rect -4100 -1411 -3838 -1399
rect -4100 -1808 -4094 -1411
rect -3844 -1808 -3838 -1411
rect -4100 -1820 -3838 -1808
rect -3722 -1411 -3460 -1399
rect -3722 -1808 -3716 -1411
rect -3466 -1808 -3460 -1411
rect -3722 -1820 -3460 -1808
rect -3344 -1411 -3082 -1399
rect -3344 -1808 -3338 -1411
rect -3088 -1808 -3082 -1411
rect -3344 -1820 -3082 -1808
rect -2966 -1411 -2704 -1399
rect -2966 -1808 -2960 -1411
rect -2710 -1808 -2704 -1411
rect -2966 -1820 -2704 -1808
rect -2588 -1411 -2326 -1399
rect -2588 -1808 -2582 -1411
rect -2332 -1808 -2326 -1411
rect -2588 -1820 -2326 -1808
rect -2210 -1411 -1948 -1399
rect -2210 -1808 -2204 -1411
rect -1954 -1808 -1948 -1411
rect -2210 -1820 -1948 -1808
rect -1832 -1411 -1570 -1399
rect -1832 -1808 -1826 -1411
rect -1576 -1808 -1570 -1411
rect -1832 -1820 -1570 -1808
rect -1454 -1411 -1192 -1399
rect -1454 -1808 -1448 -1411
rect -1198 -1808 -1192 -1411
rect -1454 -1820 -1192 -1808
rect -1076 -1411 -814 -1399
rect -1076 -1808 -1070 -1411
rect -820 -1808 -814 -1411
rect -1076 -1820 -814 -1808
rect -698 -1411 -436 -1399
rect -698 -1808 -692 -1411
rect -442 -1808 -436 -1411
rect -698 -1820 -436 -1808
rect -320 -1411 -58 -1399
rect -320 -1808 -314 -1411
rect -64 -1808 -58 -1411
rect -320 -1820 -58 -1808
rect 58 -1411 320 -1399
rect 58 -1808 64 -1411
rect 314 -1808 320 -1411
rect 58 -1820 320 -1808
rect 436 -1411 698 -1399
rect 436 -1808 442 -1411
rect 692 -1808 698 -1411
rect 436 -1820 698 -1808
rect 814 -1411 1076 -1399
rect 814 -1808 820 -1411
rect 1070 -1808 1076 -1411
rect 814 -1820 1076 -1808
rect 1192 -1411 1454 -1399
rect 1192 -1808 1198 -1411
rect 1448 -1808 1454 -1411
rect 1192 -1820 1454 -1808
rect 1570 -1411 1832 -1399
rect 1570 -1808 1576 -1411
rect 1826 -1808 1832 -1411
rect 1570 -1820 1832 -1808
rect 1948 -1411 2210 -1399
rect 1948 -1808 1954 -1411
rect 2204 -1808 2210 -1411
rect 1948 -1820 2210 -1808
rect 2326 -1411 2588 -1399
rect 2326 -1808 2332 -1411
rect 2582 -1808 2588 -1411
rect 2326 -1820 2588 -1808
rect 2704 -1411 2966 -1399
rect 2704 -1808 2710 -1411
rect 2960 -1808 2966 -1411
rect 2704 -1820 2966 -1808
rect 3082 -1411 3344 -1399
rect 3082 -1808 3088 -1411
rect 3338 -1808 3344 -1411
rect 3082 -1820 3344 -1808
rect 3460 -1411 3722 -1399
rect 3460 -1808 3466 -1411
rect 3716 -1808 3722 -1411
rect 3460 -1820 3722 -1808
rect 3838 -1411 4100 -1399
rect 3838 -1808 3844 -1411
rect 4094 -1808 4100 -1411
rect 3838 -1820 4100 -1808
rect 4216 -1411 4478 -1399
rect 4216 -1808 4222 -1411
rect 4472 -1808 4478 -1411
rect 4216 -1820 4478 -1808
rect 4594 -1411 4856 -1399
rect 4594 -1808 4600 -1411
rect 4850 -1808 4856 -1411
rect 4594 -1820 4856 -1808
rect 4972 -1411 5234 -1399
rect 4972 -1808 4978 -1411
rect 5228 -1808 5234 -1411
rect 4972 -1820 5234 -1808
rect 5350 -1411 5612 -1399
rect 5350 -1808 5356 -1411
rect 5606 -1808 5612 -1411
rect 5350 -1820 5612 -1808
rect 5728 -1411 5990 -1399
rect 5728 -1808 5734 -1411
rect 5984 -1808 5990 -1411
rect 5728 -1820 5990 -1808
rect 6106 -1411 6368 -1399
rect 6106 -1808 6112 -1411
rect 6362 -1808 6368 -1411
rect 6106 -1820 6368 -1808
rect 6484 -1411 6746 -1399
rect 6484 -1808 6490 -1411
rect 6740 -1808 6746 -1411
rect 6484 -1820 6746 -1808
rect 6862 -1411 7124 -1399
rect 6862 -1808 6868 -1411
rect 7118 -1808 7124 -1411
rect 6862 -1820 7124 -1808
rect 7240 -1411 7502 -1399
rect 7240 -1808 7246 -1411
rect 7496 -1808 7502 -1411
rect 7240 -1820 7502 -1808
rect 7618 -1411 7880 -1399
rect 7618 -1808 7624 -1411
rect 7874 -1808 7880 -1411
rect 7618 -1820 7880 -1808
rect 7996 -1411 8258 -1399
rect 7996 -1808 8002 -1411
rect 8252 -1808 8258 -1411
rect 7996 -1820 8258 -1808
rect 8374 -1411 8636 -1399
rect 8374 -1808 8380 -1411
rect 8630 -1808 8636 -1411
rect 8374 -1820 8636 -1808
rect 8752 -1411 9014 -1399
rect 8752 -1808 8758 -1411
rect 9008 -1808 9014 -1411
rect 8752 -1820 9014 -1808
rect -9014 -1948 -8752 -1936
rect -9014 -2345 -9008 -1948
rect -8758 -2345 -8752 -1948
rect -9014 -2357 -8752 -2345
rect -8636 -1948 -8374 -1936
rect -8636 -2345 -8630 -1948
rect -8380 -2345 -8374 -1948
rect -8636 -2357 -8374 -2345
rect -8258 -1948 -7996 -1936
rect -8258 -2345 -8252 -1948
rect -8002 -2345 -7996 -1948
rect -8258 -2357 -7996 -2345
rect -7880 -1948 -7618 -1936
rect -7880 -2345 -7874 -1948
rect -7624 -2345 -7618 -1948
rect -7880 -2357 -7618 -2345
rect -7502 -1948 -7240 -1936
rect -7502 -2345 -7496 -1948
rect -7246 -2345 -7240 -1948
rect -7502 -2357 -7240 -2345
rect -7124 -1948 -6862 -1936
rect -7124 -2345 -7118 -1948
rect -6868 -2345 -6862 -1948
rect -7124 -2357 -6862 -2345
rect -6746 -1948 -6484 -1936
rect -6746 -2345 -6740 -1948
rect -6490 -2345 -6484 -1948
rect -6746 -2357 -6484 -2345
rect -6368 -1948 -6106 -1936
rect -6368 -2345 -6362 -1948
rect -6112 -2345 -6106 -1948
rect -6368 -2357 -6106 -2345
rect -5990 -1948 -5728 -1936
rect -5990 -2345 -5984 -1948
rect -5734 -2345 -5728 -1948
rect -5990 -2357 -5728 -2345
rect -5612 -1948 -5350 -1936
rect -5612 -2345 -5606 -1948
rect -5356 -2345 -5350 -1948
rect -5612 -2357 -5350 -2345
rect -5234 -1948 -4972 -1936
rect -5234 -2345 -5228 -1948
rect -4978 -2345 -4972 -1948
rect -5234 -2357 -4972 -2345
rect -4856 -1948 -4594 -1936
rect -4856 -2345 -4850 -1948
rect -4600 -2345 -4594 -1948
rect -4856 -2357 -4594 -2345
rect -4478 -1948 -4216 -1936
rect -4478 -2345 -4472 -1948
rect -4222 -2345 -4216 -1948
rect -4478 -2357 -4216 -2345
rect -4100 -1948 -3838 -1936
rect -4100 -2345 -4094 -1948
rect -3844 -2345 -3838 -1948
rect -4100 -2357 -3838 -2345
rect -3722 -1948 -3460 -1936
rect -3722 -2345 -3716 -1948
rect -3466 -2345 -3460 -1948
rect -3722 -2357 -3460 -2345
rect -3344 -1948 -3082 -1936
rect -3344 -2345 -3338 -1948
rect -3088 -2345 -3082 -1948
rect -3344 -2357 -3082 -2345
rect -2966 -1948 -2704 -1936
rect -2966 -2345 -2960 -1948
rect -2710 -2345 -2704 -1948
rect -2966 -2357 -2704 -2345
rect -2588 -1948 -2326 -1936
rect -2588 -2345 -2582 -1948
rect -2332 -2345 -2326 -1948
rect -2588 -2357 -2326 -2345
rect -2210 -1948 -1948 -1936
rect -2210 -2345 -2204 -1948
rect -1954 -2345 -1948 -1948
rect -2210 -2357 -1948 -2345
rect -1832 -1948 -1570 -1936
rect -1832 -2345 -1826 -1948
rect -1576 -2345 -1570 -1948
rect -1832 -2357 -1570 -2345
rect -1454 -1948 -1192 -1936
rect -1454 -2345 -1448 -1948
rect -1198 -2345 -1192 -1948
rect -1454 -2357 -1192 -2345
rect -1076 -1948 -814 -1936
rect -1076 -2345 -1070 -1948
rect -820 -2345 -814 -1948
rect -1076 -2357 -814 -2345
rect -698 -1948 -436 -1936
rect -698 -2345 -692 -1948
rect -442 -2345 -436 -1948
rect -698 -2357 -436 -2345
rect -320 -1948 -58 -1936
rect -320 -2345 -314 -1948
rect -64 -2345 -58 -1948
rect -320 -2357 -58 -2345
rect 58 -1948 320 -1936
rect 58 -2345 64 -1948
rect 314 -2345 320 -1948
rect 58 -2357 320 -2345
rect 436 -1948 698 -1936
rect 436 -2345 442 -1948
rect 692 -2345 698 -1948
rect 436 -2357 698 -2345
rect 814 -1948 1076 -1936
rect 814 -2345 820 -1948
rect 1070 -2345 1076 -1948
rect 814 -2357 1076 -2345
rect 1192 -1948 1454 -1936
rect 1192 -2345 1198 -1948
rect 1448 -2345 1454 -1948
rect 1192 -2357 1454 -2345
rect 1570 -1948 1832 -1936
rect 1570 -2345 1576 -1948
rect 1826 -2345 1832 -1948
rect 1570 -2357 1832 -2345
rect 1948 -1948 2210 -1936
rect 1948 -2345 1954 -1948
rect 2204 -2345 2210 -1948
rect 1948 -2357 2210 -2345
rect 2326 -1948 2588 -1936
rect 2326 -2345 2332 -1948
rect 2582 -2345 2588 -1948
rect 2326 -2357 2588 -2345
rect 2704 -1948 2966 -1936
rect 2704 -2345 2710 -1948
rect 2960 -2345 2966 -1948
rect 2704 -2357 2966 -2345
rect 3082 -1948 3344 -1936
rect 3082 -2345 3088 -1948
rect 3338 -2345 3344 -1948
rect 3082 -2357 3344 -2345
rect 3460 -1948 3722 -1936
rect 3460 -2345 3466 -1948
rect 3716 -2345 3722 -1948
rect 3460 -2357 3722 -2345
rect 3838 -1948 4100 -1936
rect 3838 -2345 3844 -1948
rect 4094 -2345 4100 -1948
rect 3838 -2357 4100 -2345
rect 4216 -1948 4478 -1936
rect 4216 -2345 4222 -1948
rect 4472 -2345 4478 -1948
rect 4216 -2357 4478 -2345
rect 4594 -1948 4856 -1936
rect 4594 -2345 4600 -1948
rect 4850 -2345 4856 -1948
rect 4594 -2357 4856 -2345
rect 4972 -1948 5234 -1936
rect 4972 -2345 4978 -1948
rect 5228 -2345 5234 -1948
rect 4972 -2357 5234 -2345
rect 5350 -1948 5612 -1936
rect 5350 -2345 5356 -1948
rect 5606 -2345 5612 -1948
rect 5350 -2357 5612 -2345
rect 5728 -1948 5990 -1936
rect 5728 -2345 5734 -1948
rect 5984 -2345 5990 -1948
rect 5728 -2357 5990 -2345
rect 6106 -1948 6368 -1936
rect 6106 -2345 6112 -1948
rect 6362 -2345 6368 -1948
rect 6106 -2357 6368 -2345
rect 6484 -1948 6746 -1936
rect 6484 -2345 6490 -1948
rect 6740 -2345 6746 -1948
rect 6484 -2357 6746 -2345
rect 6862 -1948 7124 -1936
rect 6862 -2345 6868 -1948
rect 7118 -2345 7124 -1948
rect 6862 -2357 7124 -2345
rect 7240 -1948 7502 -1936
rect 7240 -2345 7246 -1948
rect 7496 -2345 7502 -1948
rect 7240 -2357 7502 -2345
rect 7618 -1948 7880 -1936
rect 7618 -2345 7624 -1948
rect 7874 -2345 7880 -1948
rect 7618 -2357 7880 -2345
rect 7996 -1948 8258 -1936
rect 7996 -2345 8002 -1948
rect 8252 -2345 8258 -1948
rect 7996 -2357 8258 -2345
rect 8374 -1948 8636 -1936
rect 8374 -2345 8380 -1948
rect 8630 -2345 8636 -1948
rect 8374 -2357 8636 -2345
rect 8752 -1948 9014 -1936
rect 8752 -2345 8758 -1948
rect 9008 -2345 9014 -1948
rect 8752 -2357 9014 -2345
rect -9014 -5167 -8752 -5155
rect -9014 -5564 -9008 -5167
rect -8758 -5564 -8752 -5167
rect -9014 -5576 -8752 -5564
rect -8636 -5167 -8374 -5155
rect -8636 -5564 -8630 -5167
rect -8380 -5564 -8374 -5167
rect -8636 -5576 -8374 -5564
rect -8258 -5167 -7996 -5155
rect -8258 -5564 -8252 -5167
rect -8002 -5564 -7996 -5167
rect -8258 -5576 -7996 -5564
rect -7880 -5167 -7618 -5155
rect -7880 -5564 -7874 -5167
rect -7624 -5564 -7618 -5167
rect -7880 -5576 -7618 -5564
rect -7502 -5167 -7240 -5155
rect -7502 -5564 -7496 -5167
rect -7246 -5564 -7240 -5167
rect -7502 -5576 -7240 -5564
rect -7124 -5167 -6862 -5155
rect -7124 -5564 -7118 -5167
rect -6868 -5564 -6862 -5167
rect -7124 -5576 -6862 -5564
rect -6746 -5167 -6484 -5155
rect -6746 -5564 -6740 -5167
rect -6490 -5564 -6484 -5167
rect -6746 -5576 -6484 -5564
rect -6368 -5167 -6106 -5155
rect -6368 -5564 -6362 -5167
rect -6112 -5564 -6106 -5167
rect -6368 -5576 -6106 -5564
rect -5990 -5167 -5728 -5155
rect -5990 -5564 -5984 -5167
rect -5734 -5564 -5728 -5167
rect -5990 -5576 -5728 -5564
rect -5612 -5167 -5350 -5155
rect -5612 -5564 -5606 -5167
rect -5356 -5564 -5350 -5167
rect -5612 -5576 -5350 -5564
rect -5234 -5167 -4972 -5155
rect -5234 -5564 -5228 -5167
rect -4978 -5564 -4972 -5167
rect -5234 -5576 -4972 -5564
rect -4856 -5167 -4594 -5155
rect -4856 -5564 -4850 -5167
rect -4600 -5564 -4594 -5167
rect -4856 -5576 -4594 -5564
rect -4478 -5167 -4216 -5155
rect -4478 -5564 -4472 -5167
rect -4222 -5564 -4216 -5167
rect -4478 -5576 -4216 -5564
rect -4100 -5167 -3838 -5155
rect -4100 -5564 -4094 -5167
rect -3844 -5564 -3838 -5167
rect -4100 -5576 -3838 -5564
rect -3722 -5167 -3460 -5155
rect -3722 -5564 -3716 -5167
rect -3466 -5564 -3460 -5167
rect -3722 -5576 -3460 -5564
rect -3344 -5167 -3082 -5155
rect -3344 -5564 -3338 -5167
rect -3088 -5564 -3082 -5167
rect -3344 -5576 -3082 -5564
rect -2966 -5167 -2704 -5155
rect -2966 -5564 -2960 -5167
rect -2710 -5564 -2704 -5167
rect -2966 -5576 -2704 -5564
rect -2588 -5167 -2326 -5155
rect -2588 -5564 -2582 -5167
rect -2332 -5564 -2326 -5167
rect -2588 -5576 -2326 -5564
rect -2210 -5167 -1948 -5155
rect -2210 -5564 -2204 -5167
rect -1954 -5564 -1948 -5167
rect -2210 -5576 -1948 -5564
rect -1832 -5167 -1570 -5155
rect -1832 -5564 -1826 -5167
rect -1576 -5564 -1570 -5167
rect -1832 -5576 -1570 -5564
rect -1454 -5167 -1192 -5155
rect -1454 -5564 -1448 -5167
rect -1198 -5564 -1192 -5167
rect -1454 -5576 -1192 -5564
rect -1076 -5167 -814 -5155
rect -1076 -5564 -1070 -5167
rect -820 -5564 -814 -5167
rect -1076 -5576 -814 -5564
rect -698 -5167 -436 -5155
rect -698 -5564 -692 -5167
rect -442 -5564 -436 -5167
rect -698 -5576 -436 -5564
rect -320 -5167 -58 -5155
rect -320 -5564 -314 -5167
rect -64 -5564 -58 -5167
rect -320 -5576 -58 -5564
rect 58 -5167 320 -5155
rect 58 -5564 64 -5167
rect 314 -5564 320 -5167
rect 58 -5576 320 -5564
rect 436 -5167 698 -5155
rect 436 -5564 442 -5167
rect 692 -5564 698 -5167
rect 436 -5576 698 -5564
rect 814 -5167 1076 -5155
rect 814 -5564 820 -5167
rect 1070 -5564 1076 -5167
rect 814 -5576 1076 -5564
rect 1192 -5167 1454 -5155
rect 1192 -5564 1198 -5167
rect 1448 -5564 1454 -5167
rect 1192 -5576 1454 -5564
rect 1570 -5167 1832 -5155
rect 1570 -5564 1576 -5167
rect 1826 -5564 1832 -5167
rect 1570 -5576 1832 -5564
rect 1948 -5167 2210 -5155
rect 1948 -5564 1954 -5167
rect 2204 -5564 2210 -5167
rect 1948 -5576 2210 -5564
rect 2326 -5167 2588 -5155
rect 2326 -5564 2332 -5167
rect 2582 -5564 2588 -5167
rect 2326 -5576 2588 -5564
rect 2704 -5167 2966 -5155
rect 2704 -5564 2710 -5167
rect 2960 -5564 2966 -5167
rect 2704 -5576 2966 -5564
rect 3082 -5167 3344 -5155
rect 3082 -5564 3088 -5167
rect 3338 -5564 3344 -5167
rect 3082 -5576 3344 -5564
rect 3460 -5167 3722 -5155
rect 3460 -5564 3466 -5167
rect 3716 -5564 3722 -5167
rect 3460 -5576 3722 -5564
rect 3838 -5167 4100 -5155
rect 3838 -5564 3844 -5167
rect 4094 -5564 4100 -5167
rect 3838 -5576 4100 -5564
rect 4216 -5167 4478 -5155
rect 4216 -5564 4222 -5167
rect 4472 -5564 4478 -5167
rect 4216 -5576 4478 -5564
rect 4594 -5167 4856 -5155
rect 4594 -5564 4600 -5167
rect 4850 -5564 4856 -5167
rect 4594 -5576 4856 -5564
rect 4972 -5167 5234 -5155
rect 4972 -5564 4978 -5167
rect 5228 -5564 5234 -5167
rect 4972 -5576 5234 -5564
rect 5350 -5167 5612 -5155
rect 5350 -5564 5356 -5167
rect 5606 -5564 5612 -5167
rect 5350 -5576 5612 -5564
rect 5728 -5167 5990 -5155
rect 5728 -5564 5734 -5167
rect 5984 -5564 5990 -5167
rect 5728 -5576 5990 -5564
rect 6106 -5167 6368 -5155
rect 6106 -5564 6112 -5167
rect 6362 -5564 6368 -5167
rect 6106 -5576 6368 -5564
rect 6484 -5167 6746 -5155
rect 6484 -5564 6490 -5167
rect 6740 -5564 6746 -5167
rect 6484 -5576 6746 -5564
rect 6862 -5167 7124 -5155
rect 6862 -5564 6868 -5167
rect 7118 -5564 7124 -5167
rect 6862 -5576 7124 -5564
rect 7240 -5167 7502 -5155
rect 7240 -5564 7246 -5167
rect 7496 -5564 7502 -5167
rect 7240 -5576 7502 -5564
rect 7618 -5167 7880 -5155
rect 7618 -5564 7624 -5167
rect 7874 -5564 7880 -5167
rect 7618 -5576 7880 -5564
rect 7996 -5167 8258 -5155
rect 7996 -5564 8002 -5167
rect 8252 -5564 8258 -5167
rect 7996 -5576 8258 -5564
rect 8374 -5167 8636 -5155
rect 8374 -5564 8380 -5167
rect 8630 -5564 8636 -5167
rect 8374 -5576 8636 -5564
rect 8752 -5167 9014 -5155
rect 8752 -5564 8758 -5167
rect 9008 -5564 9014 -5167
rect 8752 -5576 9014 -5564
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_1p41
string library sky130
string parameters w 1.410 l 14.10 m 3 nx 48 wmin 1.410 lmin 0.50 rho 2000 val 20.266k dummy 0 dw 0.0 term 188.2 sterm 0.0 caplen 0 wmax 1.410 guard 0 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} snake 0 full_metal 1 n_guard 0 hv_guard 0 vias 1 viagb 0 viagt 0 viagl 0 viagr 0
<< end >>

** sch_path: /home/vblabs/Analog/circuitos/comparador/xschem/Comparador_completo_modificado.sch
**.subckt Comparador_completo_modificado VDD VDD Vout VIN VIN VDD18 VDD18
*.ipin VDD
*.ipin VDD
*.iopin Vout
*.ipin VIN
*.ipin VIN
*.ipin VDD18
*.ipin VDD18
V1 net4 GND 1
V2 VDD GND 5
VIN VIN GND DC 0 PWL (1m 0 2m 5 3m 0)
I0 VDD net5 100n
XM3 net6 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=Lp1 W=Wp1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM9 net1 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=Lp2 W=Wp2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM13 net2 net1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=Lph W=Wph nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=Lph W=Wph nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net2 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=Lp2 W=Wp2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net7 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=Lpout W=Wpout nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM11 net7 net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=Lnout W=Wnout nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM12 net2 net4 net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=Ln1 W=Wn1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 net5 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=Ln1 W=Wn1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM1 net1 VIN net3 GND sky130_fd_pr__nfet_g5v0d10v5 L=Ln1 W=Wn1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 net6 net6 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=Ln1 W=Wn1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 net5 net5 GND GND sky130_fd_pr__nfet_g5v0d10v5 L=Ln1 W=Wn1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V3 VDD18 GND 1.8
XM10 Vout net7 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM14 Vout net7 VDD18 VDD18 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
**** begin user architecture code

.param Wn1 = 5 Ln1 = 1
.param Wp1 = 5 Lp1 = 1
.param Wp2 = 2 Lp2 = 2
.param Wph = 10 Lph = 1
.param Wnout = 10 Lnout = 1
.param Wpout = 15 Lpout = 1
.param ptemp = -40


.temp {ptemp}
.tran 100n 3.2m 1.1m

.control
foreach var1 -40 25 85
	echo temperature $var1
	alterparam ptemp =$var1
	reset
	run
	*dc Vin 0 2 0.1
	save all
	*plot vout vs vin
	meas tran rth find vin when vin=vout CROSS = 1
	meas tran rtl find vin when vin=vout CROSS = 4
	let vhist = 'rth-rtl'
	print vhist
end
.endc


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice ff

**** end user architecture code
**.ends
.GLOBAL GND
.end

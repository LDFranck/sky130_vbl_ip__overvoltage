magic
tech sky130A
magscale 1 2
timestamp 1713151348
<< error_s >>
rect 4675 4904 4685 4929
<< nwell >>
rect -18218 17203 -2751 17489
rect -18218 -3716 -17932 17203
rect -3037 14033 -2751 17203
rect 7842 14053 24078 14339
rect -3037 13747 6011 14033
rect 5725 9115 6011 13747
rect 7842 10246 8128 14053
rect 7842 9960 11647 10246
rect 5725 8829 10262 9115
rect 9976 -3716 10262 8829
rect 11361 -130 11647 9960
rect 23792 -130 24078 14053
rect 11361 -416 24078 -130
rect -18218 -4002 10262 -3716
<< nsubdiff >>
rect -18182 17433 -2831 17453
rect -18182 17399 -18100 17433
rect -2910 17399 -2831 17433
rect -18182 17379 -2831 17399
rect -18182 17373 -18108 17379
rect -18182 -3883 -18162 17373
rect -18128 -3883 -18108 17373
rect -2905 17358 -2831 17379
rect -2905 14008 -2885 17358
rect -2851 14008 -2831 17358
rect -2905 13997 -2831 14008
rect 7927 14283 24011 14303
rect 7927 14249 8003 14283
rect 23934 14249 24011 14283
rect 7927 14229 24011 14249
rect 7927 14223 8001 14229
rect -2905 13977 5975 13997
rect -2905 13943 -2831 13977
rect 5895 13943 5975 13977
rect -2905 13923 5975 13943
rect 5901 13919 5975 13923
rect 5901 9087 5921 13919
rect 5955 9087 5975 13919
rect 7927 10076 7947 14223
rect 7981 10076 8001 14223
rect 7927 10070 8001 10076
rect 23937 14223 24011 14229
rect 7927 10050 11472 10070
rect 7927 10016 8004 10050
rect 11396 10016 11472 10050
rect 7927 9996 11472 10016
rect 5901 9079 5975 9087
rect 11398 9990 11472 9996
rect 5901 9059 10225 9079
rect 5901 9025 5976 9059
rect 10148 9025 10225 9059
rect 5901 9005 10225 9025
rect -18182 -3891 -18108 -3883
rect 10151 8999 10225 9005
rect 10151 -3885 10171 8999
rect 10205 -3885 10225 8999
rect 11398 -299 11418 9990
rect 11452 -299 11472 9990
rect 11398 -305 11472 -299
rect 23937 -297 23957 14223
rect 23991 -297 24011 14223
rect 23937 -305 24011 -297
rect 11398 -325 24011 -305
rect 11398 -359 11478 -325
rect 23937 -359 24011 -325
rect 11398 -379 24011 -359
rect 10151 -3891 10225 -3885
rect -18182 -3912 10225 -3891
rect -18182 -3946 -18108 -3912
rect 10145 -3946 10225 -3912
rect -18182 -3965 10225 -3946
rect -18182 -3966 10217 -3965
<< nsubdiffcont >>
rect -18100 17399 -2910 17433
rect -18162 -3883 -18128 17373
rect -2885 14008 -2851 17358
rect 8003 14249 23934 14283
rect -2831 13943 5895 13977
rect 5921 9087 5955 13919
rect 7947 10076 7981 14223
rect 8004 10016 11396 10050
rect 5976 9025 10148 9059
rect 10171 -3885 10205 8999
rect 11418 -299 11452 9990
rect 23957 -297 23991 14223
rect 11478 -359 23937 -325
rect -18108 -3946 10145 -3912
<< locali >>
rect -18162 17399 -18100 17433
rect -2910 17399 -2851 17433
rect -18162 17373 -18128 17399
rect -2885 17358 -2851 17399
rect -2885 13977 -2851 14008
rect 7947 14249 8003 14283
rect 23934 14249 23991 14283
rect 7947 14223 7981 14249
rect -2885 13943 -2831 13977
rect 5895 13943 5955 13977
rect 5921 13919 5955 13943
rect 7947 10050 7981 10076
rect 23957 14223 23991 14249
rect 7947 10016 8004 10050
rect 11396 10016 11452 10050
rect 5921 9059 5955 9087
rect 11418 9990 11452 10016
rect 5921 9025 5976 9059
rect 10148 9025 10205 9059
rect -18162 -3912 -18128 -3883
rect 10171 8999 10205 9025
rect 11418 -325 11452 -299
rect 23957 -325 23991 -297
rect 11418 -359 11478 -325
rect 23937 -359 23991 -325
rect 10171 -3912 10205 -3885
rect -18162 -3946 -18108 -3912
rect 10145 -3945 10205 -3912
rect 10145 -3946 10204 -3945
<< metal1 >>
rect -448 9664 -438 9804
rect -381 9664 -371 9804
rect 1230 8849 1240 8989
rect 1297 8849 1307 8989
rect 4547 4901 4685 4904
rect 1227 4017 1237 4157
rect 1294 4017 1304 4157
rect 4547 1590 4674 4901
rect 4535 1533 4545 1590
rect 4685 1533 4695 1590
<< via1 >>
rect -438 9664 -381 9804
rect 1240 8849 1297 8989
rect 1237 4017 1294 4157
rect 4545 1533 4685 1590
<< metal2 >>
rect -438 9804 -381 9814
rect -381 9765 7502 9775
rect -381 9708 7362 9765
rect -381 9698 7502 9708
rect -438 9654 -381 9664
rect -438 9337 -381 9347
rect -381 9298 7292 9308
rect -381 9241 7142 9298
rect 7282 9241 7292 9298
rect -381 9231 7292 9241
rect -438 9187 -381 9197
rect 1240 8989 1297 8999
rect 1297 8951 7071 8961
rect 1297 8894 6920 8951
rect 7060 8894 7071 8951
rect 1297 8884 7071 8894
rect 1240 8839 1297 8849
rect 1240 8541 1297 8551
rect 1230 8433 1240 8510
rect 1297 8500 6847 8510
rect 1297 8443 6697 8500
rect 6837 8443 6847 8500
rect 1297 8433 6847 8443
rect 1240 8391 1297 8401
rect 7352 8170 7882 8173
rect 7352 8163 7892 8170
rect 7352 8106 7362 8163
rect 7502 8106 7892 8163
rect 7352 8099 7892 8106
rect 7352 8096 7882 8099
rect 7131 7563 7882 7569
rect 7131 7556 7934 7563
rect 7131 7499 7142 7556
rect 7282 7499 7934 7556
rect 7131 7497 7934 7499
rect 7131 7492 7882 7497
rect 6910 5974 7882 5981
rect 6910 5971 7903 5974
rect 6910 5914 6920 5971
rect 7060 5914 7903 5971
rect 6910 5904 7903 5914
rect 6686 5372 7882 5377
rect 6686 5367 7969 5372
rect 6686 5310 6697 5367
rect 6837 5310 7969 5367
rect 6686 5305 7969 5310
rect 6686 5300 7882 5305
rect 1237 4157 1294 4166
rect 1377 4141 7362 4142
rect 1294 4131 7362 4141
rect 1294 4121 7512 4131
rect 1294 4065 7362 4121
rect 1294 4064 1377 4065
rect 7502 4064 7512 4121
rect 7362 4054 7512 4064
rect 1237 4008 1294 4017
rect 7352 3783 7882 3789
rect 7352 3779 7939 3783
rect 1237 3713 1294 3723
rect 7352 3722 7362 3779
rect 7502 3722 7939 3779
rect 7352 3721 7939 3722
rect 7352 3713 7882 3721
rect 1227 3603 1237 3680
rect 7362 3712 7502 3713
rect 7576 3712 7882 3713
rect 1294 3670 7292 3680
rect 1294 3613 7142 3670
rect 7282 3613 7292 3670
rect 1294 3603 7292 3613
rect 1237 3563 1294 3573
rect 7132 3181 7882 3185
rect 7132 3175 7903 3181
rect 7132 3118 7142 3175
rect 7282 3118 7903 3175
rect 7132 3108 7903 3118
rect 4537 1597 4674 1600
rect 4537 1590 7886 1597
rect 4537 1533 4545 1590
rect 4685 1533 7919 1590
rect 4537 1527 7919 1533
rect 4537 1523 7886 1527
rect 4537 636 7882 638
rect 4537 629 7898 636
rect 4537 572 4546 629
rect 4686 597 7898 629
rect 4686 572 8482 597
rect 4537 566 8482 572
<< via2 >>
rect 7362 9708 7502 9765
rect -438 9197 -381 9337
rect 7142 9241 7282 9298
rect 6920 8894 7060 8951
rect 1240 8401 1297 8541
rect 6697 8443 6837 8500
rect 7362 8106 7502 8163
rect 7142 7499 7282 7556
rect 6920 5914 7060 5971
rect 6697 5310 6837 5367
rect 7362 4064 7502 4121
rect 7362 3722 7502 3779
rect 1237 3573 1294 3713
rect 7142 3613 7282 3670
rect 7142 3118 7282 3175
rect 4546 572 4686 629
<< metal3 >>
rect 7352 9765 7512 9775
rect 7352 9708 7362 9765
rect 7502 9708 7512 9765
rect -448 9337 -371 9342
rect -448 9197 -438 9337
rect -381 9197 -371 9337
rect -448 9192 -371 9197
rect 7131 9298 7292 9308
rect 7131 9241 7142 9298
rect 7282 9241 7292 9298
rect 6910 8951 7071 8961
rect 6910 8894 6920 8951
rect 7060 8894 7071 8951
rect 1230 8541 1307 8546
rect 1230 8401 1240 8541
rect 1297 8401 1307 8541
rect 1230 8396 1307 8401
rect 6686 8500 6847 8510
rect 6686 8443 6697 8500
rect 6837 8443 6847 8500
rect 6686 5367 6847 8443
rect 6910 5971 7071 8894
rect 7131 7556 7292 9241
rect 7352 8163 7512 9708
rect 7352 8106 7362 8163
rect 7502 8106 7512 8163
rect 7352 8096 7512 8106
rect 7131 7499 7142 7556
rect 7282 7499 7292 7556
rect 7131 7492 7292 7499
rect 6910 5914 6920 5971
rect 7060 5914 7071 5971
rect 6910 5904 7071 5914
rect 6686 5310 6697 5367
rect 6837 5310 6847 5367
rect 6686 5300 6847 5310
rect 4537 4901 4685 4974
rect 1227 3713 1304 3718
rect 1227 3573 1237 3713
rect 1294 3573 1304 3713
rect 1227 3568 1304 3573
rect 4537 1590 4674 4901
rect 7352 4121 7512 4131
rect 7352 4064 7362 4121
rect 7502 4064 7512 4121
rect 7352 3779 7512 4064
rect 7352 3722 7362 3779
rect 7502 3722 7512 3779
rect 7352 3713 7512 3722
rect 7132 3670 7292 3680
rect 7132 3613 7142 3670
rect 7282 3613 7292 3670
rect 7132 3175 7292 3613
rect 7132 3118 7142 3175
rect 7282 3118 7292 3175
rect 7132 3108 7292 3118
rect 4537 638 4685 1590
rect 4537 629 4691 638
rect 4537 572 4546 629
rect 4686 572 4691 629
rect 4537 566 4691 572
use comp_hyst  comp_hyst_0
timestamp 1713115829
transform 1 0 6716 0 1 11234
box 1667 -5363 16947 2564
use level_shifter  level_shifter_0
timestamp 1713121837
transform 1 0 6519 0 1 8816
box 1105 -2314 6378 -340
use level_shifter  level_shifter_1
timestamp 1713121837
transform 1 0 6519 0 1 6624
box 1105 -2314 6378 -340
use level_shifter  level_shifter_2
timestamp 1713121837
transform 1 0 6519 0 1 4432
box 1105 -2314 6378 -340
use level_shifter  level_shifter_4
timestamp 1713121837
transform 1 0 6519 0 1 2240
box 1105 -2314 6378 -340
use multiplexer  multiplexer_0
timestamp 1713137003
transform 1 0 -1955 0 1 209
box -199 -135 8108 13095
use vd2mux_conn  vd2mux_conn_1
timestamp 1713130350
transform 1 0 478 0 1 1
box -3578 973 -2488 12383
use voltage_divider  voltage_divider_0
timestamp 1713115829
transform 1 0 -16053 0 1 -2158
box -1259 -1438 14153 19128
<< end >>

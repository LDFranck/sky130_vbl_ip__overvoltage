magic
tech sky130A
magscale 1 2
timestamp 1713215965
<< locali >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 2319 -509 3279 -340
rect 5236 -369 6339 -340
rect 5236 -492 5457 -369
rect 6302 -492 6339 -369
rect 5236 -538 6339 -492
rect 5236 -1104 5419 -538
rect 5235 -1740 5419 -1226
rect 1183 -2314 2143 -1781
rect 5552 -2034 6339 -1774
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 5235 -2121 6339 -2034
rect 5235 -2244 5277 -2121
rect 6277 -2244 6339 -2121
rect 5235 -2314 6339 -2244
<< viali >>
rect 1223 -493 2106 -370
rect 5457 -492 6302 -369
rect 2357 -2286 3240 -2163
rect 5277 -2244 6277 -2121
<< metal1 >>
rect 1183 -370 2143 -340
rect 1183 -493 1223 -370
rect 2106 -493 2143 -370
rect 1183 -539 2143 -493
rect 5419 -369 6339 -340
rect 5419 -492 5457 -369
rect 6302 -492 6339 -369
rect 5419 -538 6339 -492
rect 1183 -758 1325 -539
rect 1353 -710 1363 -658
rect 1963 -710 1973 -658
rect 2489 -670 2499 -618
rect 3099 -670 3109 -618
rect 1183 -959 1357 -758
rect 1969 -830 2494 -746
rect 1969 -887 2205 -830
rect 2345 -887 2494 -830
rect 1969 -958 2494 -887
rect 1183 -1362 1325 -959
rect 1353 -1058 1363 -1006
rect 1963 -1058 1973 -1006
rect 2489 -1167 2505 -1151
rect 3095 -1167 3105 -1151
rect 2489 -1219 2499 -1167
rect 3099 -1219 3105 -1167
rect 1353 -1314 1363 -1262
rect 1963 -1314 1973 -1262
rect 1183 -1562 1357 -1362
rect 1969 -1427 2461 -1362
rect 1969 -1484 1985 -1427
rect 2125 -1484 2461 -1427
rect 2489 -1457 2499 -1405
rect 3099 -1457 3105 -1405
rect 2489 -1473 2504 -1457
rect 3095 -1473 3105 -1457
rect 1969 -1562 2461 -1484
rect 2462 -1562 2493 -1505
rect 1353 -1662 1363 -1610
rect 1963 -1662 1973 -1610
rect 2271 -1905 2493 -1562
rect 2489 -1953 3109 -1937
rect 2489 -2005 2499 -1953
rect 3099 -2005 3109 -1953
rect 3137 -2115 3279 -718
rect 5419 -721 5541 -538
rect 5569 -673 5579 -621
rect 6179 -673 6189 -621
rect 5419 -921 5573 -721
rect 6185 -921 6339 -721
rect 5569 -1021 5579 -969
rect 6179 -1021 6186 -969
rect 6214 -1104 6339 -921
rect 5453 -1225 6339 -1104
rect 5453 -1226 6305 -1225
rect 5453 -1400 5544 -1226
rect 5572 -1352 5578 -1300
rect 6179 -1352 6189 -1300
rect 5572 -1368 6189 -1352
rect 5453 -1599 5521 -1400
rect 5573 -1599 5583 -1400
rect 5453 -1600 5572 -1599
rect 6185 -1600 6339 -1400
rect 5569 -1700 5579 -1648
rect 6180 -1700 6190 -1648
rect 5328 -1926 5337 -1848
rect 5477 -1926 5487 -1848
rect 6218 -2034 6339 -1600
rect 2319 -2163 3279 -2115
rect 2319 -2286 2357 -2163
rect 3240 -2286 3279 -2163
rect 2319 -2314 3279 -2286
rect 5235 -2121 6339 -2034
rect 5235 -2244 5277 -2121
rect 6277 -2244 6339 -2121
rect 5235 -2314 6339 -2244
<< via1 >>
rect 1363 -710 1963 -658
rect 2499 -670 3099 -618
rect 2205 -887 2345 -830
rect 1363 -1058 1963 -1006
rect 2499 -1219 3099 -1167
rect 1363 -1314 1963 -1262
rect 1985 -1484 2125 -1427
rect 2499 -1457 3099 -1405
rect 1363 -1662 1963 -1610
rect 2499 -2005 3099 -1953
rect 5579 -673 6179 -621
rect 5579 -1021 6179 -969
rect 5578 -1352 6179 -1300
rect 5521 -1599 5573 -1400
rect 5579 -1700 6180 -1648
rect 5337 -1926 5477 -1848
<< metal2 >>
rect 2499 -616 6179 -606
rect 2499 -618 5340 -616
rect 1363 -657 2135 -643
rect 1363 -658 1985 -657
rect 1963 -710 1985 -658
rect 1363 -714 1985 -710
rect 2125 -714 2135 -657
rect 3099 -670 5340 -618
rect 2499 -673 5340 -670
rect 5480 -621 6179 -616
rect 5480 -673 5579 -621
rect 2499 -683 6179 -673
rect 1363 -720 2135 -714
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -897 2355 -887
rect 5328 -969 6179 -959
rect 1363 -1006 2135 -996
rect 1963 -1058 1985 -1006
rect 1363 -1063 1985 -1058
rect 2125 -1063 2135 -1006
rect 5328 -1026 5338 -969
rect 5478 -1021 5579 -969
rect 5478 -1026 6179 -1021
rect 5328 -1036 6179 -1026
rect 1363 -1068 2135 -1063
rect 1363 -1073 2125 -1068
rect 2499 -1164 5488 -1157
rect 2499 -1167 5338 -1164
rect 3099 -1219 5338 -1167
rect 2499 -1221 5338 -1219
rect 5478 -1221 5488 -1164
rect 2499 -1229 5488 -1221
rect 1363 -1257 2355 -1247
rect 1363 -1262 2205 -1257
rect 1963 -1314 2205 -1262
rect 2345 -1314 2355 -1257
rect 1363 -1324 2355 -1314
rect 5328 -1294 6179 -1285
rect 5328 -1351 5338 -1294
rect 5478 -1300 6179 -1294
rect 5478 -1351 5578 -1300
rect 5328 -1352 5578 -1351
rect 5328 -1362 6179 -1352
rect 2499 -1400 5573 -1390
rect 2499 -1405 3177 -1400
rect 1975 -1427 2135 -1417
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 3099 -1457 3177 -1405
rect 3317 -1457 5521 -1400
rect 2499 -1467 5521 -1457
rect 1975 -1494 2135 -1484
rect 1363 -1610 2355 -1600
rect 5521 -1609 5573 -1599
rect 1963 -1662 2205 -1610
rect 1363 -1667 2205 -1662
rect 2345 -1667 2355 -1610
rect 1363 -1672 2355 -1667
rect 5328 -1648 6180 -1638
rect 5328 -1705 5338 -1648
rect 5478 -1700 5579 -1648
rect 5478 -1705 6180 -1700
rect 5328 -1715 6180 -1705
rect 5337 -1848 5477 -1838
rect 5337 -1936 5477 -1926
rect 2499 -1952 3327 -1943
rect 2499 -1953 3177 -1952
rect 3099 -2005 3177 -1953
rect 2499 -2009 3177 -2005
rect 3317 -2009 3327 -1952
rect 2499 -2015 3327 -2009
<< via2 >>
rect 1985 -714 2125 -657
rect 5340 -673 5480 -616
rect 2205 -887 2345 -830
rect 1985 -1063 2125 -1006
rect 5338 -1026 5478 -969
rect 5338 -1221 5478 -1164
rect 2205 -1314 2345 -1257
rect 5338 -1351 5478 -1294
rect 1985 -1484 2125 -1427
rect 3177 -1457 3317 -1400
rect 2205 -1667 2345 -1610
rect 5338 -1705 5478 -1648
rect 5337 -1926 5477 -1848
rect 3177 -2009 3317 -1952
<< metal3 >>
rect 5328 -616 5489 -606
rect 1975 -657 2135 -648
rect 1975 -714 1985 -657
rect 2125 -714 2135 -657
rect 1975 -1006 2135 -714
rect 5328 -673 5340 -616
rect 5480 -673 5489 -616
rect 1975 -1063 1985 -1006
rect 2125 -1063 2135 -1006
rect 1975 -1427 2135 -1063
rect 1975 -1484 1985 -1427
rect 2125 -1484 2135 -1427
rect 1975 -1494 2135 -1484
rect 2195 -830 2355 -820
rect 2195 -887 2205 -830
rect 2345 -887 2355 -830
rect 2195 -1257 2355 -887
rect 2195 -1314 2205 -1257
rect 2345 -1314 2355 -1257
rect 2195 -1610 2355 -1314
rect 5328 -969 5489 -673
rect 5328 -1026 5338 -969
rect 5478 -1026 5489 -969
rect 5328 -1164 5489 -1026
rect 5328 -1221 5338 -1164
rect 5478 -1221 5489 -1164
rect 5328 -1294 5489 -1221
rect 5328 -1351 5338 -1294
rect 5478 -1351 5489 -1294
rect 2195 -1667 2205 -1610
rect 2345 -1667 2355 -1610
rect 2195 -1672 2355 -1667
rect 3167 -1400 3327 -1390
rect 3167 -1457 3177 -1400
rect 3317 -1457 3327 -1400
rect 3167 -1952 3327 -1457
rect 3167 -2009 3177 -1952
rect 3317 -2009 3327 -1952
rect 3167 -2014 3327 -2009
rect 5328 -1648 5489 -1351
rect 5328 -1705 5338 -1648
rect 5478 -1705 5489 -1648
rect 5328 -1848 5489 -1705
rect 5328 -1926 5337 -1848
rect 5477 -1926 5489 -1848
rect 5328 -2015 5489 -1926
use sky130_fd_pr__diode_pw2nd_05v5_37RBXE  sky130_fd_pr__diode_pw2nd_05v5_37RBXE_0
timestamp 1713020003
transform 0 1 5406 -1 0 -1887
box -183 -208 183 208
use sky130_fd_pr__nfet_01v8_MG6U6H  sky130_fd_pr__nfet_01v8_MG6U6H_0
timestamp 1713020003
transform 1 0 5878 0 1 -1500
box -496 -310 496 310
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_0
timestamp 1713020003
transform -1 0 2799 0 1 -1705
box -528 -458 528 458
use sky130_fd_pr__nfet_g5v0d10v5_EEVBR7  sky130_fd_pr__nfet_g5v0d10v5_EEVBR7_1
timestamp 1713020003
transform -1 0 2799 0 1 -919
box -528 -458 528 458
use sky130_fd_pr__pfet_01v8_J2L9Q3  sky130_fd_pr__pfet_01v8_J2L9Q3_0
timestamp 1713020003
transform 1 0 5878 0 1 -821
box -496 -319 496 319
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_0
timestamp 1713020003
transform 1 0 1663 0 -1 -1462
box -558 -397 558 397
use sky130_fd_pr__pfet_g5v0d10v5_YHAZV5  sky130_fd_pr__pfet_g5v0d10v5_YHAZV5_1
timestamp 1713020003
transform 1 0 1663 0 -1 -858
box -558 -397 558 397
<< labels >>
flabel space 1105 -1255 2221 -461 0 FreeSans 1600 0 0 0 M3
flabel space 2271 -1377 3327 -461 0 FreeSans 1600 0 0 0 M5
flabel space 2271 -2163 3327 -1247 0 FreeSans 1600 0 0 0 M6
flabel metal1 1183 -539 2143 -340 0 FreeSans 1600 0 0 0 avdd
port 1 nsew
flabel metal2 1363 -1662 1963 -1610 0 FreeSans 800 0 0 0 out_b
port 2 nsew
flabel metal2 1363 -710 1963 -658 0 FreeSans 800 0 0 0 out
port 3 nsew
flabel space 1105 -1859 2221 -1065 0 FreeSans 1600 0 0 0 M4
flabel metal2 3317 -1467 3773 -1390 0 FreeSans 800 0 0 0 in_b
flabel metal1 2319 -2314 3279 -2115 0 FreeSans 1600 0 0 0 avss
port 4 nsew
flabel space 5419 -538 6379 -340 0 FreeSans 1600 0 0 0 dvdd
port 5 nsew
flabel metal3 5328 -2015 5489 -1926 0 FreeSans 1600 0 0 0 in
port 6 nsew
flabel space 5383 -1810 6375 -1190 0 FreeSans 1600 0 0 0 M1
flabel space 5383 -1140 6375 -502 0 FreeSans 1600 0 0 0 M2
flabel metal1 5235 -2313 6339 -2244 0 FreeSans 1600 0 0 0 dvss
port 7 nsew
<< end >>
